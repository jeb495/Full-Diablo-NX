MPQ    6�    h�  h                                                                                 &8I=qH
�_�c���n�t�0Њ�������]nɬi����^Ƅ,���ě(�X~�y��q���ܕ)B�`~�Y~/='�(�H�t�:��Q1���c��8�p3�$Ҝ��0��B3�8���:���MW�8<���]�l���)�p��13�����6S(��O�b~x��5%9�%�����H���~�2t"Cur
S�����hyǿi�������X���w7���`����5�.��n/Y�&d^��r��a��nLe+-���kWV��)�+���B�jnZ�:��zd����L�-J(ub��T��k^�r� s�|��!���xX^��Z㎬6t�y�p�6!�H�쀛�@J�:�_�%n.J�l)����ԎF. �y�.��-�$��"��:��X|��o�E�K��C	Xc�0b2;��=�����R,�Y@���h���N�#7G�����D/n��%i
�Q5��m�<{�P���	;N��OTj_�G�U�#B,�rM�0�W�s
�Fe��"�Yx�>hJ���0�~�.�@��x�k�d�1�ާz�={�t�<���x�)���E6���d������%�,Аv���}N�J''���q9�S�F��16h�@�w���zV���Yo���/羴�bUV�R��LV�:�ه
��0x.9�BD�1zN�X>����J���"�����U���K�rJ?m���	���Dc��`w�.�����c��4�����%X�p4�$/c��M@�i��@���a�QF�&j�ܳZ���� 4��*��b'̐^m����rE$k������T(n��74���fJ;�Il�V��f�g������~�b���ā���\T�Zy�2rI���1#q�O�j�a���X��+�hC� jjZ���w���d�]��F�M�]�*��/fo.O�>�=J|ġ��3�V�^��_A��m�
4�A2�/ Jt~@������[�M��/�h��@0�|B��!
z�}q�����d�$��z�x�w��s|�G.���T������.�٥a�6}������
�|7"�radEs	W��3!����@x�e%�W�6�ͬ�ic(�x�=i����y�P�]1��$2��m��,8�u��C`�k�9u�U9d��*��� %���"�<�*q/*�k���Z��L:|h�!]���w�?YBAQ��P@7����Nf�b(	M,��������k��~�#\�d���wWB-�[������h��$'�y������ Ã2�+��T��&.�ʹ��}�~]G}(�.y���(>I(z +�8sr�)��R�^�z�˘\4�*�,5���`%|t��	钸擪oK��'����|�E
�u���ܺ�3�P�a��U}N�DK ���~��W���T�LK�y����|vY���!"�О�X���Q0ݦ]xlIij0��̯a�L�l� ���#���xH��zS3-(�r�J���jx�V_1����@�#DZ"��dN\�����L�f�z�� �s�0��D�}Bp4�Z}��K���ĸk�Ⱥ�y�x�a�Pe��R�E�r�X&��3��.C���Mδ��C���ĥW�~U&gf�d����6>�gsq�i����Y�Dw؋�2�`Ut@{g6��C w ��cP{�*(���*�ݕ�:ync����/�����l`H��5Q�/���y<S`�_����Iv�re\x������G�I
��L��?�����j^�(mʧ �q�QTõX�Q��V`ݯ�"W�v#�8L�뫺�=-��֔ �ɾ�l��~�W��!=Å=�M5̌�ʿ���]e$ԼC@`��_��B% � g����d� �`�#�I)�tv8�*�7�N�t���_�G0+�T\����x�F� D�4mƫy�����?�qz �?t���U"������Z����L��h�۰(����.e�v��x{��ώ"�L&'��J�[ܲⷄ10��j��r
&���y�����Y��|^Ptz���[Z�ԇQ��i����p�z�X�r���m�ظ�=�ܴ��G��f.D���#��YCG3y���ɒ^
ќZ�{�R]5vk�Z��)���BTS0xRW�j�
?�m��
��{{��ʱ����H`��Bb���v>�Sp���w>B���.#`��4��yg���6Pet�̣r�N�r8�����΍,P�,*�LBy��[�w��S?�R����`�½8p�:�8�����#��{^�f�Ųvp5���ʦr?D���xL�R����&KibY���u�1Un����(\Q~�OdQ!+�Bz7�{8��~l����ő�a�^p�!� ��dj_H�bƻ�g�W�ݯ$4W~|]����.p1�KMqE��a��64��|4OWx'JX߰XR��S�1X��Ș꧎+��lr9=!�H�Q�ƭ2^�� 1��<���H�0�B��`&T��,�J[A	��A%K�r�v����.��aetU�z��p�ۺ��*ݯ�W��=��¯Ǹu�Ʀ��v �73���#6�������k5��K����
sԗ^,7TY�ֆ��j��,�猓�Ȋ�lp�Z��bH=צ]���5<���U员����˟M�Ln� /��k�v�qq��LK@Cν����n����U�����jI��r���d���b^��zϊ6�x���w����ڔڢ4��tEp/a.r�2t%����n�����Na�j�/������Zw#(�FY5���j�0i�^;=�����_�<�Hv:&�R��%��-Q�P�Kc~6���p᜷H���J����<���7�>&��)�� ������e&O�8��T\�j��0�6��wi�qK�аٯ��4*] l���_1��;z᷊��H3�E A?"������qb��w�s� w��@�X2T�d��'d��F�4��P�J��VA�~b]���V˾���!0u�D�� 7�~s�b�. ���Ճ��N�}��I���X�(��\��n��b0�o2�QuU��B��ɟH�D�d�1��	�.d�5�ě�+­V,�
�� �`�뉄�:���rs�҆�k�HG�!vS�0�!����F{���t{F@��2l!�T�3�=<���ŷ��d�r 	���5ǚ��7���e�]Ԙ�i�Ý��I�Xz�}����`]�MO�!0RK�,a�b���_�hSC�P��x]~��p��-k���|�ɣI�9ct=ީr�Qo��ۓ̣��`~���A�W��%���8 ���5Ƨ�ѩ�A�A_^�"��P�/�)��+HT�j V�P�f����8�nU J��_�[�8L�H4J}Gb�Pb��&�ݽsݡp�R�i�D\0Xy>vZ^��O���F�6���Gp��$U�<_��.%fldv�Ė��F)ۦy9IW���7$�"}Xz:���|G�qox{K	�����X�S�06&�2��x�c�`���n�t�0��ئFX(h���i�#7�����Dj�[�W.��Q�Nm�C��k�*������T�K�G7�3#=�r��0P����
3�����Y��h�؝�+��~M q@������zi�ނ�zx}Xt �����l)��E�\����Ҕ+J����,��Xh��x�J_n���^���u�} ��!9h1q�f@^���.V\`X�ދ�v�9�/�=}��gL�;���e�V)3w��]fO�������y5�����Ӽ��"� �{�Ƹ�׺��3m��	74���Ζ[�0.s���jc�����J� -�̫x�$��<�ȌS��.��|*ׄ₡�̊[�>��hϱ�R�*���s���j�yy��eT�E���M��g�#n�n,���Ȍf;AE�х�f�HZ��-��!	~���;d\���\o��Z��.r$�B�l���	t�\j�ҳ�^��@�h^�j���z0��b����F�QR޸�֠��,J�o�
Q>�hW|�'�ԓ��V�_���a��(��4J2$6�JOTL��P+�6[���Y�hy6�@K_fBm��������蠑��_+2���x��i��uG��+y$�T5_X����.�;�aA�H}��W�$6
\d�"�IKd�%.Wt��3к�i��@3�@��h�͇��i��x2�e����qPP�@���^�q]X�[I,sK��}��.u9��U����E	������<��/�ɛ�%ZP�u�t��<md��k�ܸA���P�� ��#�f]��(��ݛ0�l�`[�F�2��\~u!���g��-fj�����i����*��+o���K2?�����A�G�4��}���|�(�զ�r>�!j �(s�G��X\��9�-��u4�]d�'�i�v�+.���ؒ3qx�J���Y�X�~�F�w
6�Ȑ��Nc��x}UX��k, E�~~���l�K���X��v4i�\>�c֎S���Ձ�a��ld�j��h��f������n���;�4ؚ�j�xc1�z�	�-D�Ʌ�����VZ���I��A��#_��`��N7�Z���;��f���[�����D)�kB�oZ������R�X|k���;�JxL�-P�$RD�������w�ΣM.>ɋƨJ?�{K�����Wpa�&B��d L~��)�>�Aq8�}V1�.AS��2[=Bt{�g�,KC꧒J6�P6�Z(�k�*���p�y�汈���*֞��`��f�P/�^S�T8�<����IѮ�e����7'��ܗ
���LAS?R� �qja�((� ��̭	�3pQǙ�`x۱��vv~�8/��g�VA�o4Qnl+�i�R9!�lp=�"u̧���:�X�8D�$w��a	�Z�,B�ԩ "n�njڛ�1��6B)�9�8Y�l�7�N�s�Y��br���Ὦ�$_�b�Dd�ƦD��f�lcR ���Dn��5q���k��nD�7��#�'�C6]�s�}e�_�BKЎ_c&t�	�ֶ[��f���4�����d��>Q����=���|y>kzB�\�6;.��Mo�.�����r��-y����S��=�ht�P���2��f)���$��pO3�{�7Y^�@`��
���mvf@��V;��<�Tn�)R�x�j����0���N�{vF��Z�?�'`�LSb;�6�ޱ����+�->=�m։�`�~�9[�gw�&6+��t+��>~N�`������',k",*j:BTⷄ��-wN��S:�s�K��`Y��8*�?:+ܲ�yj���G�,�(Y1® �Bp�%���L?���nM�Lɦ���>&F��Y���uZ+�p��
9���\�݉O���+��z�$a8{b�6#(q�l5ka"�p5���|�2����Hjr���Ȅ���$o�`|�������1�5M,���|�eڱi����4�׭'��=�+�R᯹�Wy����"-�g��9x�HFDUƨx�^f� �G�W��ft��
���Ta4,�El,	���%�e����aEe�<KH�^��x9۵��*8���l�X2*�*)�ujW�g� _k8�܂�68��u�k���Ƥ{�fF��Ҿ,��9�����������b��d��@��
\�Ag���r��Ω�Mm��HQ�:�Mu�J�;Н��<v�b�x��>yC�v�.(.n�6ج��hK���e��������dӷ�b�]�z�ry��s!��$��x�����R}JpJ��rRV�%�)~��}:Ш;oN\\��A&��h��@w��WF4s/�V���ˉ�^o��X ��}"< ?W:���Rmx��1%��t�cy5��l�Qp�FH�s|Jr������~��$&�[0�Q*v�C ��1.O����A\$���T��6��:i3�`���l5��qB�*8�l�ܸ_̄�;uAъ�x�H�@7 \�Y"�o
��k-q�Ҁ���1�� �X����Af'��%�!0�4����8�Q�AZ4�]���qC��H]j`�D%v7��y4�bb�� HJ������pۭ�I#�XS���WwMn��60�懣l�Y�T�Τ��ؠ>d~M�qi��l5��Ķ��(���q�[Z>���넦�:���(?Ѝ�^�5��#��!�Ź0��׮��QF֔�Y��{aO�׭^�/=低<�о�ob�p�۫*�0e�ܔ�ȷj��\;��{Ø/�x+�FL�2b�ATu]^���F���E��'�����Q�S^}��ELD~�ݲ��A���ږ�����NV��QtX��r pC�����ޫ޿�0���g��gX��������f}5�@���w��E}�^��k��^ ��ߥ+c�6��
V]ZF��Q��x�?nPz��E�9��jL�ĢJ��b�?`�,�ᗨ��s��G­�)����X���Z�O��������6�h΢����p_�0�. K�l�V��1�F$�&y��ҕ@$JB"�8:���|��Fo���KE��T�KX�dS0QN�21Ľ�>SK�8ެ��-�m���Jh��!ۄ�+7=W��G�D��ݜ�V� ��Q�	mrjc����������%T�WVG�\�#8�rj�0Vxq�
�?彙:bYh�כ�&s�~�1�@r���i�����]����t����n)J�E�$����5��w��,Fˢ�<��s��J����8���Z��)���1��@��-��arV���\���Ʃ������yL�����c��m��!�x�B�'a)��ߏ����ӷ��"y��6�����j�h�4mg��	r��zD�V�.��$�M�6c��|���u`����$e�N����m��74z��å�G���1 �)��LGx�Tx�?�g��0퐔�͒��EڈQ�?�y���n�c�<_�G��;(X��L�hf��]����EN~��I��#W͉�2\��nZo�r�w�#ܧ��5�W����䐂vhy��j`[�U�ڹ�+ȓɐF��3���Id�e��o$�>y��|:���.��VÀ`��E���4�2�\bJ*J�-;kƩ�[������h4�@fxB�e���+5���Ѡ,�Z�{�B�2xS�멎uG�Tp�Tp&�N�.Ͻ�a��;}E�����
�k="]@%d��FW��3Q���Y@�[��x�r�b3�i��|x�&���Ȏy�PeC���������6a�,�3��
��9+WU�_}�`^��c���<Q�/`$���Z�L���r�W����K��~�Aǀ�Pv�;�ٜ9f���(t�KW���/�!�\����8½-!���ƶ�^3���y�2��_���O2��,�y�S�\�ʯ��}�����('���L6>�:: �F�s�#9�ӻT�?��A͂4"��"_j�`L�����wP���%�F����w2�r}x
�4m�Kr��i��Wn�U3B�񺫄 �+�~ySnNs��QPK�/��8v\%���Z3�N�"��H�Sl�j'��xa��B<���h���y�Ȓ�%�ux~�`z��-����H�ؠiVUI���<��-P#z�*��N���Zn�Ktf�(p��AJ����DD�Bf�nZ���ߏ�a�k��z��<�x{IP�5�R����5ۡ�
9�im?.9ƶ��Ɉ6s����cW�c�&�d[�O�l^�>�תqm�ڍ8	-9���26:_t�,�gl̚C}뒥(@P���(�`�*$,�K��y�4�:Ϫ%b��j �`x���k�Z/B��/��<ɜؔ��&.rI,��e��"��h�=�
��mL|�?��e�j�$�(�g �G'|��Q^�`'���/vٱ`8���#��J��?=*l�>��Mí!�5;=t����ʵ�L�C$JQ�v���UBB��i ݏ,�!���5����J)(�8�G�W�NP�7���}���J���myu�R�D��ơ/���,����55ﺎ5���� x�$o�8���װ^n���e���Ve��Ɏ�u&�<l�m�m[��zE�����Bu@w��
�јs^��	$|�L�z��]�<I��i�ǟ���)��0iİ�:ۈ��|��є=�ً�}���f$�!�UF��ϼ;3�_���x�^˗ߜ�<\�0va�]�w��ŉ�T��cRM+cj����mڟ@3�{q���g�׈��S`�b��j�����Z���>8���G��9�CT �g�-n6�tfA����#N�n�^Q��K��,��*�B/�Ä�6�w��S5z���Ʉ`��8EF�:��9�TF�F ���T�9�{ٮp��� SO?:�0I�0LϤ2��&A'YM�uEU������ʷZ\�\+O��k+��z�&86��G?���G�a]�'pФ��w�\��4H%�@���)�	_�C%$�aW|��}����1D�@M�Iܗ b�,�+�l��4�w'Sy���AR<�_`�����ꝯ��B�%9�W�H�Vƣ��^�� �P�rn���_̾�d=�W�sT��#�@�	CN\%�9ݴ�zi��{"�Q����"�۰��*�����s��¥�GuE4J ��u��I�6p���0X�k7g��Aq��A����,m�r�̊B�I�h���}�����{��Gl���n�ܐ!���J�ʉ���L���!��p�MP�7�v� �uv�U'�H��P�Cru���n��Z�˳6�G�`��X�Ռ��d��bTV�z�z��v��]���6��X(���pe�br͙4%cܜ��/�CNW�Q���Ȩ\�_�&/w%F�T���x�f��^���o+'�~�<U`:��RH�ÔV��� -ctTȲ��pW?H�t[J�C�}���Z7��t+�&�E���S6��tz��O��X��\\_�]6�=yi��u�xo,Pg���*�l2"�_gqa;p���>�CH��L wz"u%ՠ �q�WĀ�[4��|I�{u�X�Л˚��'�?���!45;݌���LA�	�]zc���������j�D`s?7P�tWb�� ��j��DWE��H�I^�eX�9��R#�nR�0Z}���1����C�A�Kd������5�0��I�£/+��}���A&���:D��d��Шۡ�|�V���!�Wu07^���:F1A�1{|~(�(q/�
���+�<� ��G��H��n��J���9���ğ���9�'Ó��-s�Γb�Mg謁�U]9����g5�`ǆ"=��)�Symү�?~�@����cV��t�Y��寵Otst+r{�#�����uȿ:!���k'�i���@��������5|��L/����^��B�Ѹ�Yl+~�̇`�VV8���0.��.nK}�����ѝ�L�`yJs&/b�NN�gʑ�C �s�K���逺[�X�,�ZTnr�A��ŝ4�A_�6�����{�q:k���_�.ۯ�l�Vr�̋�F�by�ݍ���@$5�="s9|:|�=|��ooT=8K�
7��s�X<�50l�"2�����s�^���"�������hKd۟�;7�����D�	������<QF�m-�����h�z�T��Gm�#3A
r^p70�'�1z�
l�t��Y)�h���!e�~cA@-o糼]�p8��8Oy��,tVy��O�)�TKEg���3Ҋ�1���,���1��n�lJ]�X����o��sO�ג1��@�6�����V����^[�/^���,o�w�L'���ʁW��h������y�������8Ӳr�"�ѐ��4����AmB{M	���Y�Q3 .)�`���c�����莶���!a$ ߘ��j.�z����]�%��s���E	�d�����������f���S���
�[��E�G�zaR𝙃n�x�H���Ɓ;C���ǚxf��p�G8����~�����r�D��\��Z�u+rڌԴ��ߧ Y��R���i���=̊h��j�n0��P���.�)F���n+O�E���Ko���>T�|u����|�V��ŉpS��s�4:��2�%J`�ha�0[�<�@P�h��@�۱Bc�f����.�o��tIU���=sx�T��G�Gc]/��T�T��.�_�a�a} ���L�
R�b"8W�d��SW�1�3�c�չ@�$~v}�-��=��i�	xh�&�䉎Կ P f��3�g�1��M,�;������9���UjU�{������r
�<��/���~�Z��kƍ�r��G��A�A��P�N��5�fJ
(:8͛fHI�Vxi���}/��\��	��x���-�籼(�Ӻ��ҵy*�T�����2��r�4�[�w�*�?}kj��(�B���F�>Zt� \��s���N;x��d�|�4�`A�$�黰�V뭔�^P�)�� ���P�ߴs��m|
�����Ġ�眢҃�U��� {�~t����C؅W8K(Q�N�v��1������͎I��b�o�ׯVl��j��тS|F�}���[�����
���x�7z��^-�������;:VP����ԛ#�t�V*QN�}[�0�T��&,f}�*��U�a�D_� B�y�Z�D�3�?���
k}^���x�7IP���R:lul���	��W�.4�]�^�T��b�	"�Wf�j&�[�d��5�� >���qȿ����L,c�It2W�t��g��C0� ;6P�F�(�u�*��r�&��yM���Y �"��=�`3�Zӆ�/~E��
�<kp�0%��v6I�_�e�s� ��YX
|�L���?��F�yj�F(�f� �������GQ=B;`�����$v4p�8}"��{�����%��z,'laG�Hm�!N�=/,��ݺ��0¬��a$�K��c�P��B6�) �/��<|ڑ�x���c)c$�8�����zN����{��V���L-�H���b�D�jƜ:'���ٝM��a械E<�iU��Z�c����u]Bؙ9�yƭ�iA�e�w���cx����&*�N�(N�[-����a�sl�}������v9��^=�`�|�z�z8|���\�8��:v#��`�����t��
2�I�=b�c����h�f�����a��)3�cf�- *^�O����#�Fv\������D_T��%R��bjw�����7{lV���,u��p�`�lb1��E}��IT�ar�>3j��?
"����o�Qgm��6�l�t��P�t��NȜO��>�9,�b�*`b�B
@���w�_�S0s���`���8`�v:!���/�8�J�L�b��O�ͮ��pfc���y?��$L?�B����&<��Y���u�~��aS BI�۫\��O5��+�N=zH7�8�������>�"��a�:zpk���r�uW�H����6W45�n��$�b|.M����B1�~kM�u�ܲ2ڧ4V�G#W4 8�'�@1ЁPR��E��!���p��|�9�"�H|��ƞd^R� bA-��v��\k��������T�O�;��	���%|�ش�mԲW����v�)��*۫��*�!�L"��Ν� L�u ��L � �2��0�6ˤ{���ikR0|Ǽ]��
�H��,���<��ޫ�]���ފ�=��n.��u�w���LM�i��|0�gz�0�@M+b4�ʷ��)�v�����}�WC��$��n��8����["���v��GpZd	��b�n�z`��)�]�H��{�ڳ�����p�!�rH�v%>�+������NR���@�����q%w���F�N
�����+�^�6���έ9�<6��:��LR#��G��!��co�&�"
�p�(H��JhO�XX�����b<&�OR��ր��#��)vO�2]qh\�H ���C6�4i�n��3o�k^�g��*�.lm�k_~�;ka؊���Hd6� �\�"����{�Tq��H�(���̖�?�Xc�˵�7'�U&���4p�!�ޒGMhA�F]5짓��>�����D��|7�5�ob�� �;>�&@��]����I�wX��>�M�n�2�04������)�Z�IN�d�<���~�?g�5?r���º�̜ڛ�pш�ܫ��zJr:�����>��?M���n��k !'
%0�W�����F���j�{��ף��� �3��<Ui��?n�u?QQj�9����S�~�����w�Î��.P	Љ��h���7�]u0��:6#����sh���"VS�}�;S�~xÅ�!������z'7ɴ��j9t�oxr��iL�T^F��1盪���č;���6��O���5W���Z@4�{T�^��U�a�A�Z��+�g���}�VB��0�쮌unFΠ�������zL��J�eEb\},���5��q�s��j�c�urX���Z��!�6� ����6C��X�[�,uU�#�_���.�4qlw!�g��F�ZyJX�����$P$"�Y�:W��|���o��ZK��
X��{0��22'{���p��*��E��]��Wih@�ۺIT73��a3NDK��(���\Q���m����D���QZ��TVдG�##.��r��m0��L�'
����O�!Yd?Sh�4��w0~^�y@��)��q<������)D�t�"h��,�) рE"��1���sw�d-�,��)F��i.�Jp>��Z��H!��o1"�@/�z��'[Vmw��Ë�3���7�δ�>��L��ſ~g�+d���F�ȴ�w%�*��Q��ӭ{"/����1���^�ZmY�	蟊��ÖL�.�J=��F`c)(>�rP���g)�\�$�
��	���I�����3���=嚒y�ܟW�ςT˫�-����N����]����5E�&���8��n�d��4Ƚ%G;^� �B�f\�������{�~��c�L���nD\�W�Ze�+r������0�Mk���ݰ��AVh��XjV��p~���C��.�F����ɀ��E��o��>/�|�z��d*�V�"'�˂�Y��4U��2�	�J��Ќ��\���[�= ����h�@��Bި��Ͱ�i���b��P�ö�tx�>p�� MG�_�
h�T���U�.�!�aRc�}����h
���"��d1�TWE��3�z@d���n�K�טiOݪx���<�/	Pۨ��,�/� ��Z,$d��NB��7�9�;2U%�p�Hq�$�MB�<�7A/�9=y��Za�2&��]���Х�$�A=�XP��Y���fn"�(����C��6���{j h\Og����hx�]-�V	�C2�T&�ҐJ(eH��]���>2P%y��z'Ȓ2Qʥ0�}FN�3:m(]����`�>��z 0Ns�;������<�ܷ�y4X�	��5��s��eؒ��n��>��
�d�O�һh�
Gsx������[�M�PU��<�0�� �~o)u�T�@}dKC.ɧ��v�[����iۍ�D������ݒ`�l�{oj���.�6ĸH���hE����E	����x���z���-���6k���ډVK�N�Zde�r��#��ыMN��k���ZfxV!�l.!�>Dz�B\&RZ�Kќnht�)�kx���L3x}-P��	R�c�G��Do���`�./ �ƹ߈�"I�$�BW�ȉ&��d�S/��'T>��Rq#ǀ��ΐG���2�)t,��g�kbC��[mlPgă(��6*u���myZ06�pD�~�� �=`�jӡ�/�h.���<?Y|���A���I��eH����3��
W(^L�ޜ?#����jrkX(Y�� #�=z���iQxF�`I���Uv�NB88��&\�� ���;�l�:�C7�!�(q=�`����ʫy�ɠ�$�e�&E�K�B�� S��W3��J��)�I8*�Ķ
��N2��x���P�@2g�#�2�2�D5S�Ɨe}�w!��sڤ���+vU�D�>����<%����X��[�T�d��>2���ebb@��C��B�&�ݱ��9g[H#�p���N�ĸ�jvH���Nj��E�@|��@z���ǝ��s���Yr������0�^ш�C/��j�==̓�w�`xf��	�E��3凬���4^����F����vW�Q�-�[��#�T��oRC��jRR�YHk�v\�{g���2�p`&�ub�� jݱ?с���>.�J֚�☯+����g�a6�jt�G4���N��d�Lם��,�2�*�5�B�J,�GS/w��S+���\u`��8{�:��k�
Ի��x-����J}}�1�gp!2��6�?0�S���Lzcj�h,�&7e�Yru�ث��{���\=��O�++���z��Q8������G���a��p���mT%��;
H�a˻��~��IWl$ �|������k1���M]p�̈́R�"�,�"h 4;�'�(?�\R��kֈu�<�`�P���k9)>H��ƙ

^w�� R����U�ז ��z���y�T2��6_�	�Nw%7QX��G��H��ͼ$A6�IS�ۦ�,*Iݭ�2���̓�u��=�,� 0Ƙ��7;6&������km��7j�����ԃ��,�������������~��
�����Nq�Dh���g�#J�AD�&[���9MTA���b�P��v	t�NY�8��C:�l����nZ��Ao扆VU@�	 �Nd$bJ�sz;�"�d����
�vT�j���W�p��7rÀ�%�*�Zv�yNMW)曚��ҙ��#w��F��O�1�ܜ��^��f�%2����<Q��:��R��!���ه���cj���}H�p��H ��J�f��3LH���H���L&�ym�bW�t~���U�O�6x8d\��o�%w�6�kiD���u���'*�g\l�c_���;f!Ɗ�VoH�� �^�"�_�V�0qNXE��j���r�1*�X��ШL'������4�Q����>B��Ak�]�ķ��k�깏����D֟.7���j7�bs- y�~�AЉ�:�=���I��X$˚�H�}n�s0�
a��mW��H<�5c��u�dO����5s���5�Ӆ�\%�Z�v��PwZ��u�_:�c>�ڎ����`�r��b%!b��0mqɮ�J�F������{�<���m����n��<�톾�W���V~T@�T�/��T��Y>��I�[�og�Éx�����D�[������{]�l���-���ՆY��#�K;S�������~Sf��\����u����~�%�Lt���rq��DST̏gX�pb:���}�Q�� Q�0����b52�\ѕT���|^������r��E+�XЇV��V��	�RO��I�nA� �V�
�GYL�^Ji��b7�����͗y�bs�u�¾7j�0�:X��ZJ�]}�;���w��6��γm\���c�ղ_��.��lP����Fy��ĕqjZ$k��"i��:2A�|3�o��UK����eހX�V&0��+2���㫁�����.��Y�h�;��ռt7�z<�WDV�ܜÐ��T�Q���m�����{G�p��5JT�<rG�׎#)�`r�c0<+ig��
%`�*�9Y��jhQ����~�%�@��P��6f���|8d��t��D��)\)[m�E�;{�L��ҀuI�?�,�|�z��d�9J��]���3d��i����lg1]!L@�U�����V�i[�NB�)a�%o}��\�y��L]������ޚ���&������Rx�e.���0Ө�'"�B�g?���U���m�VS	#Y�K�E�G�.߽��~%kcDޤ���7�l̗�a$6Vզ����0��h��NGc���U�m�K��&?������P�(�	�͐�齒Q��Ek%d�����Ӽ�n������x�;y]���/=f70Ȥ��W���~��ڱ�!ͺy\۹WZ��r�'�X���V(˃HV'�(����eh�'[j��9�oH�ƏM�d��F�i �$�G�zf��>�o�8�>
T�|�!����V����&#���4p�2��J����4��[������heQ9@�םBYz��h�����Ǡ���K���S
5x� P��%Gu|���T!<����.��a��T}v=��H
HB�"��Sdl.JW�e3����Mz@�M��>�r���حi�`x�tH������1P���G�S]����,_������z9<�U�������O6�(�:<�/1��t��Z�T�����=�Nu��'�Ax;pPG�\���|f�P(�͛�F�LƲ��i�\��R��+��t-R��^����O��k������Y����2�s?𪔷ȭ��� ��}!R�n��(�ﵦ���>G� ���s�w]�D����[��c4����U�q���*>���ۃ���9�E[���̆�c�W
�B.�|B����¢��U���k,� ��p~j�_������K^+B�D�~v�;�H+&�%�?Z]����M1�l�c�jw��	�����S�'����Y{�V9pxϽ�zx#c-o���q,'�q��VFݳ��i�-�#���LvN����_>��DfsT��Ԭ�א>D���B��5Zd�.��?}��=�ks9��PAx8�P��R0{}"��Q6�:��.*} �|j�g�3�? ~W\+5&���dA=�=�>��q~i��b�?��2���tg�.g=k�C�����P"b�( �*�d��t�y�3���@<��{"`���ӼQ�/t�O��C*<zg��f���h�I=��e���6$[�VI
2��L-��?����j�>
(�� >���Sܵ��;Q�j�`��?�	��v�LS8�6�A]��(���C��j�l�"��>!�!R�=��]�s��&����$��G���F�jB�e� π�r
�ڇ��j��)َp8�rg�w�Na�E���κ~߻7M��7��m�DЪ ƒ�����ZOi��������:�����D��������A��֞�_X�e=m38��A��	#�&�ݔ�E�[cȷ�q��)����hs����ѩ��� nE|�6�z.�h����Ԯ~��p]���.�A��@���t�?�=ؓ�<��ΪfN��fj�� cY3 �Z�#o�^\\����S�Y] vR����Gź[1T��AR�j-�!���џ��{b�N�x��+ֱ`A�&b'I�v=�zy����7>)������jy���gc�6���t�k̪�%N�XV�oy��|ʼ,�";*V))B�����w�J�S&�Ϣ�r�`Eu�8�w�:���Ή�A�����E�I���p� ��QEG?�'�p�L�7F��G&24�Y^��uFR}ܣ��*[��\x�Ok��+�bz�ɷ8g�:����ذ.a��p��^�h�Æ+@uHV�%J���$($[�|dfj���01U�!M�P���Fڝ�����4v�'$0�W�RMY��.��WZ��Q,��{�9d�H�NƔ��^�<� ؂������R���w5~���T����1�	T��%�\���²Mߢʨ"9|#��䛐ۡ;�*�����xh�����hu��[�X� �y~��^�6����am)k�",ǲ����uԾ��,>�-�� ]�Z!���o�s���8�[��S`׭�?���0�*��+�9Ě&X�M�e^�'E"���Ov��8���H�CUpd���n5j�|\��E?�Q���i��սKd?�Hb���zR���@�~]�q0��iG�>�Gp�A~r>$�%�����v��R�NH@��������_*h*w��nF��%�B�d�7L4^�~7��e���8�<lWl:���R�[ٔ��~�W�#ceq��ئjp�-IH;8�J^�I�`\��ߨE/�&��侽���/3#��^O*�O\]Ӵ�Xy6�i�����΄��]�*�њl�n_8�;aP�O65Hګe ȀU"�E�1�<q�Ԁ~":����4FX�q���)'��W��o/4���Q�=�A�I]�����cO�4��wK�DfT7!1�exsb΍� 4�B�\�����˭\*I�VX���C�pnc)�0�G��;��	�z�$��Q�d����D���5�U��"��ed�Qa+G7)�pn�:UE�������g���ㅏy!��`0�_����FB�Ezj{�ˎיh_���1���<��������+��v:�oXn��ò4�_���
w{Ä{������<>��6@�-��]ʄ��2A4Yp��'Y)c��t>S���1�~.)����4��p9��jp���t��*r�)����ʐ������7S�z4��qo�K�7�uL�5��ЈZ౫�^��/��c�ІX+�i>���Vɩ@������n<�����e�lL!�mJ�D�b;��IZ�uxs�:~��*���X �;Z�m%X/��v=���16C���|��J�ܧ4_y��.l��l�ĝb�Fby �@�,pM$�~�"��y:��|n~�o%U(K�*���RXm�40�.2���V�$�-�{�����j�h|W��O�7)q>��D�-��^9��0QW7m^E����r���[�T���G>�1#$vfroC0�\��U�
}�v��!Y�MVh���0~��@^E[����^���C��ht'֙��FN)�)�E��h�g�]�������,2��_�Y�_ފJ&������N�~��ʕh��1���@e���m4V#|�H��2>��'���$Y��`L��-λ�aj�¤��&"����-�@�������ӣ�6"���"���#q	�TA�m�t�	^2t�ߖBZ.:Q��9$c_�3�hc��Gٲ�ҭ�$��Ǧ��9ً�C�#���i��3��HA���ϸ�~��;R���~����� �3�� EFD��+��n�n�w�Y�
�3E�;��{�8��f������@�~��a��u��\�;�Z[f1rk�����#��?m�Ca�z�}�n��h�%jL�Q��b�����F�?R��Ԡ5��і�o��>�+|&�Ԛ�gV�Dމ��{��v�4�Y�2�6�J�a��@�2L\[��ܪQ�`h � @�PB�k��C�������_�F���� �x?���3EG����T\����HO.��a��}1��(��
��Z"�[�d��3W{�x3���0��@ګ�ǀkdEU����i�w)x9y=�Lv��%zPQ�8�baذ��=,�������X9��IU��t�̲�����<=�!/��6o�ZB��08�Ýx���aJ�A���P��W����f$33(kC���P��_ƍ�&��\����d
.,-���y�J�)�F��P�%uS��<�2���e�����ʛ98}�u�X�(�vʦ���>k�; ��1s�9Ͽyk�����-�@4�Ց�3F�̝��z�.Ԁ��%�� �|߅)ӻ^}/
�1�7��ҢC��U�U��� L��~el��6ض(�KyH���z�v{�7����� ��:���s�$�"�l�k�j�ڂ�g�.�ҷ���$J���s��vx갇z�y�-J��ɬ+��qVA�4�{��W#�Ǯ�N~���KA�!�fnÙ"����"D�}LBR�eZ?#\��6Z�_vkn�0�B/x�-�PFR����SȰ�ӷ.%�;�o���"R"�Z�AW׭l&�q�dGN_��p�>�7kq�5��$�}��|*2�m�t�ͻg؊
C	S�2�P�I(,u�*k�ݷ��y�V���9x	�ֵf`d��ױo/�]���<����=�lI�X�e��%�Qo��)�
�Lh1�?Yg��uhj(2\(�"l Y�*3M��z��Q�t`����kvEk$8�+�\~pmwֶJ+�l2Y(�9+�!_�'=`*�.<ʡV�~R$6��Ip�A�pBG�j ��O؍���}�E�)��8`�� |N�P9 ݃�T�6]߮���S;Dk"�ƍ^�-��
��i��!7��t�����r�b��;�n���ʻ��ʎ���e��B�`I�]�$�&;���Yqq[~�t�fx ����.���I��z����$�| ŗz��}���������ſ򜂝�ԁ׈����=�d�w���9]5f�j�����/�30q��V�^73>��E���V�vM�5����u��T�*�R95�j6L�ϢL���{]�m�Ӳ��n`\/�b���֣ͱ�Ay�2��>$S��P%�%�@��2gޏ�6r��tR���E�+N��#���u�7�%,�2�*�<�B�0U���twU��S!ݢ�e` ��8�r�:�t���r��*��3��@�1�禠p�//�l+�?&�&�I�L�+֤��&-#Y���u��tUq��6�\���O�"+�uzY��8"�?xu�%�ų�7aI�*p<+o�c>ކ�d�H�f�!�vs ����$���|�"���.�1��M��E����U���Q�4�8�'�W��r�R��xL��r���q*���M9�D�HM�'Ə��^-� �����Nd��M�Rt�C�Th��,��	�ϒ%���F�ȕ�ʃ���d�nۜ�%*����}߁��(��vu�*��b fM��å�6ܷ��_/k�K��-��Q���2�,��Ʈ��r����Z�5����آ6��ĵC�Hw����u^�
��3��T���:�M����b�����v��;�}�Ю۳CpZ��ˆnGE���wRŬ�L��čw�xi`dZ�Rb@x0z��y���.�H܋ln\��DϘ��Ap��r���%��x���Я�NCI��Q�T�H�gE9w�RF{���}C����^�R$�۸��j��<��:J]R��@��&ׇ��c`��3%�pCwHV��Jُ9��@�F4J���u&�-��9���y�!oO}�G�+\K+�[Z�6�QMi��̅d.U���&j*[�lw�_�c2;\v��5H�� �¸"�J�4yq�ؖ��V��迖�^�X��\���'�f��hO�4!���E8��A!��]f���{�ꯦ�R�9DLL�7�ތ`�b)  �~��w�5�01f�7`IJ�$XZܚ�>�n�Լ0Fѣ�)�������|�M�d�g���QP�F5p��=��a��,�@�>����k0O:�F�P���,��hZ?�j��!���0�n��D�F�2� 2�{�z��ܦvfa���<&WN��������X���T�w�|�8U���u祦���?wLк
e���@����]����mt1�
E�p������S�m���M�~	��8�Ϭ��k�f��H囄Zt� �rg���N��8��#)���D��7��,�q�f���Ua5�a��{�L��^���r���/+��LV��G����� [n7�4�L�����L<�J_�b��g�S�ڗ�&s���t 뀦��X�.Z@Xy3iy������96����i���]����^_��(.G�-lƗg�8�Fݫy[���畄$�[�"_{:�@{|�	]o�G�K�b3�ɄX(��0���2�}��9r�_���B��0�h�yh7�&��7����D����
���Q��m�����fE#�K�Tu	G�#�r�ɐ0��3���
�]ٽ�%�Yh����m�~ohc@"J�(nc\V�ޤ*��*Gt��f�ʃ�)"ES�YԂ^|�vڑ���,m�q�Cx�Z�wJ��YD��iث�_���CƇ1ӱw@ �R��@;V~��*�Ms�� m�_���C�L��ζ9xy��˿��F������~E��n�"O!ӞVB"@3r��FB�>|źϯ�m���	�+�����=CP.����Bmcz���7�"�����$lM򦪦���?��D'������#���P%#�S�\����̴��אb�GQ�E!�v�f
>�	`�n���v���;�����D2f��_�3��L�~�b��]��0��\ސZ�K6rF :������wǃ>����D�)cQh "�j�6��̹<�]Ț��F�5���@���c��o��>�	�|a��5�;V�4��É��b�4���2��Jq�e�T����E[�������h�l@�S*BO}��0��W�3C�AUr�	W�x��[�0l�GkR��yT��<�&�.�'!ac'}�6wCC
>q0"��xd��WX3�}���F;@��-� �7�ͩ<i �xԝ�����@��P1��}[�S���}��,՜:����`T9�UV]����}@��ީ�<x��/g�wjhZrOPW����m��vՂ�<��A�W�P}^K���@fk�(&�ݛ�tc�B2��h����\ y���H�n�-�b輔�ٺ���!�V���\����2ap� ($������}׹`�o(.7��n�>ƙl H~ys/P~�:y?�[��h�4)眶	x��'��B�ޔI;��PR�l����%� ���Y��
XA���̠�o���1UzZ)���K �q�~`Z� �q��K����:[vV˄���:sގ5�&��U���2Nl��jm����'��i�&��AՓݕt�VZ��Px�ezn�-%k���ا�	V<5��k6S���3#�~BpKNY���X��R�=fin�}��MԋD�f�B���Z�Y�N��Jki���]S�x�j1P"�R&
6�W̡�uN�p=. ����Ԁ���u^�WRP0&dcd�{��sE>���q4���f5�K�5j:2}
�t�}gs��C�;C�lďP��(G
�*���ݒ�;y���A��1s`����19/j�V�v	<��X������ I�@ey�0�l�%��j
��L��m?����	hj�EN(��� t,��fN�UE�Q)�`����OQv���8i��w�J�љ֑�f)dlͯ#�4U!�S=���I����f�Zy$qt}��<��B�n+ ��"ب��}ٗ� h)Oya8��u��ִN���E���߱������� D�wƈ������Ŵ�.V5���i����F[������*��a؅|&��f0�U�e��i}d���.��D�&�>����[�h)��M�߃��i�@Gr���f�_L��v�:|sz$���X "�$��Ǧį��|���t��〈*�׊5@G=�Oٲl���f2���C�v736��^�^*n����p�vH.b�> }�0+T�~R���j�׆�
�۟G� {X�(�.�,���O`w��bd,�����)C��p�>6�֫S���t��gYx�6M��t�����L
N��́%4U����,c3*Lp)Bvӑ���Ew��S��m��`���8̍F:��]��64H���3;�5�Bj-pR^T�1�?��R�B�L+@�9��&(2�Y��u��lf���<�\��O�߬+��?z��#8�))T���Ŏ.1a�#Npל��^�t��KH�p:�<�]�����$�+V|��U����1|XM� _�;(ړJ���4�x5'Z�����Rn_���t�������_9ڏVH�Ɗ�I^��� ND������Hٹ�-��~�T��'r]	
��%h��3zѲCl��^N�����cۗS�*Z�;�8f?���f��u�\�8� A��67���p�k���ǨO���M5�4�h,tJ���D;��x�I���P�����J���7��@W�{�6����r[�o#.�=lM����?��!<jv�k;�D��i��C�dL��n�C���lJ�d҆G������3��du�$b�Aź��gǯ�R��g̪�b阴Q�p���r4˹%�:�����J�N>rO�x�5�`�Ow��BFV�����;�m��^�F-�6,��%�<���:��eR��X�3�㇍Z6c[������p��yHqZ�JTTu��������{|�&���s�����<��O��ɬ�\��v��{�6���iU���)�zDS�]*ZHlY\�_n��;W!8�U!HP�� �$�"|p����q�ȍ���+���3�B��XO}w�!0<'xW��CO�4\�|���S3eBA|d]!����{�*�{-�2D�R�7W�[[Z�b��� �*X��ٗ�����xI���X�?�9_�n�Q0O��8���\|���:jd ?������5+���X��
~\��&�esH&��fQ:hX���/����E�!m0>~����F�~�	P{J&׏��Qh��X<�;���_���\�=����������z��-Q�@�K�z�����u�Ϩ�`	�#'�]�i��ǂ����	#c���|E�S �t�'�~�m���j��f�� A(�V�'t���r��:�����@C�A�ě�_R�0[���lx��c��kF5�u��FQQ��`^}����T��F��+��ǏGV��mz�gn2�ȡgż�x�LLWM�Jڣ�b�x��=O�J�s�$���ī�a
�X6��Z�bY�Z��G��HN�6��k��{��g�0_oQ=."��l8��ӑFx�y�������$�X�"�u:��R|�*o[ZVK���v�X�h~0�ޅ2i��`����C����t}a����h���&�7��͊�D����\��sQ�m��~�(VB�����)TBA�Gtr #�%r%p�0m ?��]
s*����bYPܩh"o����~�9@��C��mM�1�pt]	����)lXEsOԝ�"��<��4J,�z
��.�UJ���ȍ��B���>#�#`1�[@�����3�V� ���X�h�F���:��*G�L.��α����(P�>���	���0��y��$�ә�I"��j���O�Y���J>8m�	�D��[�8�b.����dc��ɿ^�������H�$�T���m�A����c��ꩂ)�p����܋TS������a�ʸ:M��6NW����E����D���(n���W�ȩ�;ʂ�.��f��änR����o~��豸?���Y\,�)ZQQ�r!��	% �'�ك9�
�0�J��X-h�jB^�w/��wAd�5y�F�K��5���J�po�|>��|�Sc�� V�慉7��En4�?�2��JL�b��2h]G[�-*��Th��{@�,Bʮ>����U���FR<�$�d��x���K�]G�vפT�qɬ�2.�i�a��N}��^a\
�8r"��d��W�13�����@P����]ZJ�̈́�Mi;��xo�����u���kP��[Øu��K��X�#,E'��@J�9M�aUR�������5��a-<�DS/�e��Z�|����]������9A)oP�6λ�f��y(��+��O~��p?�C�Ve�\�i���L��z-�Qм����@�:��m�Q�[��غV2��ۡ ��6Oʑ¯}�}�(�����>!s} ��sJ�*ϵ��6�Wܣj�4� �ݜ邆�y��d�I����Gf�����߻B4�T��
�pȭ2����9�~UU�-��� �y[~[UTpZ�,T�K��]��[v1�!��������0LU�)���~cFl!��j�}���XĤ��$���&��
堇x �Kz�D- m��"0��B=�V7����8�^��#��Q�N4��W�c��hfd2U�؇е��D�o�BH�Z�z'�Z����9vkd�4����xiǥP=�R��4����0�Ȱ��.T��%1����=aW��&?ugd��߼:>�'�q�$N���	�*�w�2X��t^rg*�C����v�PS�(b�8*aW��mL�yF�*�ܮo6P`�����/�6<�Q�<+R5�7����INI�e4���e���
�_ L��?�����j�x�(E@y ���)�ɵ0��Qd�`������rv�8$�a�� mV�l����lh&w�/��!�^=�s'�d��ʗ���5܏$��{�7��B�"� ?.���Oz���=��{�)��8������Nr��v�҃���,�����:D�q�ƃQ/����
��Ic}�x����\��q��h��~$$�@]/� _U���ze�M��*N������&�>��(�[�K�\妆��hĤ|�j��rVѺ���1�+|6A�z��3�]�_���A(ߣ�S��R�
�Je�Eh���=��t��S�o�Rf�7�w�l�1)|3QX֏���^�@��2
��*�vC�
��3��T+)�R/��j��ѬE}~��.#{S.�ʉk�\�T`�+b�!�]~�+2A�h�L>9f��g��"��~�gԀ�6(��t���{��N�bS������$,(��*�ËBQ�>�3�w���S0��;W`v`�8��:��a�v�h�q]y�i�6MV��MZp��W�?o�k[�Lft��Z�&#a�Yo�auw�-w�g8�ns\)�ZO<�+��fz*8���DP���i�a�mepr.��Y���<�H�`�Wz3l����$��|5����.)1f$MI���9�`@򎻆4'��'����R^(�����1����dk�9�H�f�ƅ��^�8 	�Ó�Äz�&����>T�CK�"c-	eЮ%# ��Ne��b��9�-G3��5qے�*�
V�����Sug��s�� �T����6�d�����k��P�#�g�ciH�oA�,������ku�F��kЊv�[���:���~*��v�sU��-����b/��_�Mr[��������v�S�I,��$a�C��<����n�`[�-%Q�$��Ba.�z�����d���b6�z�I�P*��O}�bJ��z�c�o:ap��r�Θ%����F�t���N9���|���{�nw�?F1���Յ��z^�ZR���r����<�y�:�\�RjV �nϤ�(�cV�����p�j8H��J�8���[y���S�&�as����`��WF�Os4��˳\�붴���6� i�����M�1���*5϶l�a
_	�+;Ra��`�GH�� �w"�5�����q:ٸ�O	����c��X
3��<�q'�g��o4��e�"+`.;�Aש�]��.��=9L�D�x~7�"V�lb�n� e�����&^���+�I��|X�m��4��nt��0��ѣ)f��zN?Ρ&u�\d��+��Q��5暨�s ��J��d�����T�a�:f�v�Ɓ��J��^I<� ~�!Ne�0�󮘾�FS�v�{9��
�|�,���Z{�<\@v�����<�������m
��ű��5�`��eH�uDL�۹�0��%����X][�?��:(*��Q2:˶�7�	S����g~�1?�H�̖a���{Y���xt7sr]�c����{�i��dx��#|ꋞ娢#�������W5��%с�����^x:�(÷��)+ ]9�B$\VZ�Ŕ>��n-P���^��3Z�Lr�JU�
b�G���緗��s�I��*�l�Z�XQ��Z6���<L�'�ʸ�6����k���z-ު_���.���l<���nY4F39y�4�]A�$�u�"Uܤ:��z|�Lo���K�Nښ�3	X�Y�0�2�tu�;����L]:x��[@h�j��A�G7�8��DBq��/���@Qh�m����C4��\h6��=T}-qG�k#��r�6�0(��P
������Y��h�M1���~%+�@�;Գ^�0R�>�ZX�P�t�Ri��])��E�IԸ|Q�l�
��,ㇷ0�}�PV&J7)���$�����UR���h1I�s@6Ѿ�F}V4s`y�苃=����<�ej%L�ά�(.�="�5�N��y�¾�Q'��X�Ӕ�M"����S��t�U���md� 	~)�H>�3�.K���j��c��п�����̃r$��裂bٜ�w�T�b�����.��\��ƣWω%!���<��>����r�QZ�=P*E�`I�ܞl�?��nזj�L�d�_;�y1���Wf�8�������~��бߵͦ�h\G�jZ�vDr���D�<��F��4B$ҋ����nMh6�5j��bR��������[{F��pސ��f)�"_0o�f3>v?�|�ٶ�kn�V��Ӊ��%� ��4���2��J'��ʓYa[��z�b4�hQl/@#PWBE ����o�ij�7c��#�xpGx�f>VGa.Q�T*�\��.��aJb}b��y��
4  "Z�^dX7�WL+�3�� �A��@S#�|��_ �ivO�x
G����ߎ��P��#ó�sI���3��,KH�U���9��MU̿����s�x��9�<�j/��`�Z(�Dͺg�n��l�@��r1Ad�VP��ζk�f5<�(�n��K��8������N�\Vz��pO?�->`\��pͺ�5��F���(���ө�2���;�����}��iZ��(d���»>|ln ���se�?�0�+����t�4_j��a�ݪ#�)��iz�EQ�"@��1��V�H�O`
�F�hm��&t𢴤xU0Db�W� ��~Vp���j��?K�_��0|�v�4zpx��+2`���;�9��l<D�jcw0�u�y��+��c��׽��]�B�x;J:zd=�-��y�]q��ݥ�V2a�!��]�#7	�8S�N����Ђ�<f_yx�3�\�×�D�B�d�Z�VŜ���0x�k_�@��9x$D�PX"R��EW�k7��p�.1wƀ���S	��<�WH�[&��d�5>��N?>�Ϣq��эUl��4+�^23�mtS֛g���C�X�"I=Pp(}��*����H��y����w�/t���Mu`����(��/`��,O�<f����F|��~I�q-e������м
�=�L�2?*I[���j9�( �� �8���p�7eQ�;`P�O��m�vV�8�����������GS�g{l�"�*	�!p7J=�H��cv�����$������2�jBX�� ����ަ��s.p��K)��81e���N��1t��:�ߧ���jKU�Yd�D<I��~2�>�J;���d����Hɺ��,���<�C2��ޝ�bF��]��wb�K+e��`�s8����&L"芴�[�N���K���z��m^}�f�ڞ�������|Q/�z�6��IԚ���ܫF��J�a� �`A[�+==�G��([U�
��f�(�үu��U�3l%�Ϳ^�w��m���v>(/��8�ŦzTF��R���j�{,���5�}�{N�s��XɈ!~`��|b��gꞱfZs���>\��a8i�V�	gO��6�.t��bON�P���n4�hm�,C#�*B7�B,y[�nJDw&��S��#�`1D8$�:P=�QY����>���1ђ��P'p��㽝�?�x.F��L�Ⱦ�o6�&��Yʼ�u2ylH���\�R�\dW�O�L�+�
�zjo8S�_l�����D,�a��pp�p�T����"HBp�r���Ҹ�8�$G�H|�����^1��M6��T��ډ�s�i� 4bY�'��N��R��}��2����?�t9P�HYaƀ(^>� ąA�/GG�>P'��`���(LT9��t�	� �%�;��i� �9y���+h�$�P��ۍ�m*f�Ӧ�0�����uB^��IX 7�F��:�6���M��k��Ǟ���>�+Ԫ�),�g������&���"������?���m�u���4O�q�,o1���
ݘ�����JMM�s����W�v�[�35��SUC��ԟgn��.�h��#F�=4����[թ��d�� b���z�1ռ�����k�]�����=�*C�p"�r*�c%`@���o�ЀhIN4$ �b?�y<��ԕwv�GF��.�cܣ^َ���rڭ��<�o:y�RE?������Q)cQ�J�D`�pt�H��WJJ=��z�͙����I�&�+[�)���F��rO�*
`\��,�6}��i����ɥI��*�5lφf_�i;M�����H�� 4I�"r�՝�Nqu	��@���	P����X�y�W*o'n�K����4�9����D)1XA2_3]�h��I�H� ���6tD��t7���Q�b:O�  �}��t��$~���I�X+���/WVnϖ[0wH�D� ��_.�|g��VdV�P�ܨ�a��5��Ď9t� �ڽPb3&~���\6i:�
u����e8����܅�P!��I0t�i���-F�w1F{9H�ׅr���Q��<�d�4񗫟�A��ۀ���G����V�p��v���pǒP����3r�
��]6$f��!Ś@����������S6~��h�~�t����9�}��\�s�֑����Mt0��r�㘊���̶u`�w5D������]�q����a2�5y�Ѽ���^sɵ��Q���-M+;�Ǉ�ؼV5�<�y�e�P�Yn(�����>L�%�JЂ�b~6�����s��vm-���dXl^8Z�׽��M�b���~'�6��M�zz@��u�H0�_e\j.��lw؂�	AF��ylְ���$� "м�:y��|Zk�o���K��w�,�[XYjX0)�2	���d����s#��y�chh[�\ܐ7�����D}r�K�@(Q�dmJ ��^2���)�|�T�9�G�y�#��r�u0�c��9)
i#ʽq��Y��MhXL�����~�<.@Jxo�y�3����5� �1�t�������)"[�E��F��;��a����,�x�ad�K��J���uN��v$���,��<�1���@�S���y�V�4c�����I϶�������Ld�Χ�x�Qhƥi�Pg����y���u���/PӏQM"Q�������]*�@��m?,�	J�8R�8�.��.�މ�%_?c�L �T	��<̾~x$=�¦�c���߳�'��L�����P,�0�$|��#������V�l����E�������Dnҋ��_��>; �ӗ$�<f~a���<��3T~�BT�n���a��\b�SZG�Mrמ?�%��]�&�/����{�Z��hQ� j8_�-O��Wm�k^�F~�2�� Ƞ!�E=7�o�A�>Q��|�~�܈V���$����/4��2w�Jy�E��[��窽��hC�@>��B�qc������+t���2>��;x+�,�זG��h,OkTH�^��Bu.�M�atV}��I�
�':"5w�d�	bW�Dx3�x���]@�ʜ3}pP���:�i�,x������Q��P=���	��f��H�,������u���9�yU�M��8]��o1�<)�/8yK[ñZ�7���?�/�t������A��PNO�α�If���(WU�#f���MP��?�W�\�/�ִ��XJ-�����v�6��Ҳ?�����#��θ�2r�`�Q��4��ʇ�W}hE&��(�Ѝ�}��>ׅ? y�s���ϫ7D��5���@4�ێ����8�9s�n��03���"��9��l%������J}�
i/��#�̠A&��/�U���-� ���~Q�,&o�آ�K��X���ov�ZL�oca+Ȏ&8G��E��$clW̬j�ЂP�
�n۷Z:�Ψ��g�V���xV�0z��-���ɘ��x.cV-�R�|(���#Rg��t�N����<V�#0XfZ�י����~��D�xB>�Z�R3��S����kZӨ�nG�x��:PsV�R��ui������A:�..���I#�1��[�W���&��'d3ð�D�>���qE�u��	���r2�t�n�gDI�C�|�};�P�V(���*Wh��#|7y�#�����E�Bk:`P�Cr/�����,<��J�m����'I��e�j��ے��w
y;�LTVs?�)���j�?�(�� ��,sD��ߧQ���`����,jv�$�8�f���B�����"��7El�s&�%�n!� =L=�̚�Yʍ�!�빍$"��Nh�-=aB��m �������.����) �a8�����N(=�~X�Ue=�"3�E���T
D�@��y���������e�9��f�L���\�ޔ���S����ض~m�6�W��A�e���.�t��g~&����E`�[�qx�R�}�p%�K�����&�pN��?�|l='z�����������wO棍a���x���30�y(�2��so���N����@��c�{��~-��I�)��mQivސ�#�f=\�$G�Ѣ���Y���}atlf�&��;]���{��R��k�*G�<�g���@e�fp��K�ox允��(��a�
-���8"p,Ś����	���S4>��50��O/RZn߱
C��z��Z=NR�E_�!�^5�g.�s�����1�:�,� �Ĉt�lw�7ZmgCDl�}��|Zu�y~�A�s<_O�tX�hjZw	�(�c�����/��AC}�������f����Q�(W0F�S�7��Y&�B����$(�ݕ���Y�FĠ Em���,���Ķ�6F�)(&�M�������T�O�c"N��<��]��5H�����v0P��G�O�h�B�|����3ԣ�ܕD��34~��1p�i�n! �`jPC��j	_��O���N�"nz�HM.��63�D�|!�(ȼ�@*N{����o����8��ݪ�6�}��AH�9g~䐧tJ1|f������'�˅㔬�]z�➨�@��狵�?"=W�GP�r�(˲ME]%{"�<b/��o.���7��l��{�Zp�O��������DB�e���7ƌ�<������n��-�_ �#*D�Q����[���<���5����~� VC�8�	8b��s���t6�j�0���9�M�5�i�i�ހu���-�̤pm�%=w/�����şq/{&����DC���q��'RU�3�R��2 X���T�����g��b�� ���R֓��kdvG����)�|R�/ɽ�&Lo�V�0��sy<��:�߬�!�Qg��>���-�Z�g}�yC���_sK�|��X��S�[�T:.��lC�a]��/�7�w`��-5P�S��_ػ�Q��&UdM�o-5�?n��;`�/ۅ}9��E/QD֍�	��#��-��#�я�2/P����TO������o��d��?�k�d-\5�6�	�\-��Y*�d�ۊl�Ԣ��]��H���Y�n�_����nVFϥu�x�s&�-���2u���V/мw�nA��Sr5�
��!�ȝyIi9
����@z5,�EC#�:�a�ov�ȃ�^���.ZY�Ź��"}�}?8���kZS��g�ufͯ�o��R�E#�"����4�b��=��|3[F��oRf�t����mhF �J�IG
h�|��!@p6����G��@N�7>seIR?���!�v&�k#p�$W�M�TQ7����ɦ�0%�_ѭ�\#�4!��!@u}
4�������>�#C0��U\-�B:�!W��`]�kTf������]��q���Y�׆��XD/���n���8��;0�r.^�Y,��܉E<)!�h��d�tq�r����/�T�	vAvU�	>ܓ�Fl<�3l���O���k������z[�7�>؏e#��P�
�os3����9�(����GM�݄�����e��֦$H����.�(��*�&����S�ţ��$e�r�*�(R79j]6ƅ�?�dg��Z\�#(W��p��G��N�L"G�mN�+?5	�D����DO��<Y�P�7YpLL����=~�R����Ɨ� ����^��n�&�jj���2��3���+*�Ch�q.׍gr �����M���2xUX�E`�8ω����'�l "�(%e�0�e4�}��Zwk�;E7�������˟p�����y��(�EEZ�n���?lу�e���AE��ZJ��W��1�מ8=N��<�B���S2 Y���F�9�%�Hc��o��5��\ƁOSf/�F��[\̧\ʴ�/���| ���?��h[l�	�T�[%a.����cl��75��v�w|h��6�{��AY�K�ª� }5��L�����f�?�ߏj���'F���f��s���ș=�?�رn�I=a۫�����霗���H�b��1���e?���vNu���{��sh.�2o�u�:���5���* v�P[T�h�;*J�FТ.�q�_��҉H�gKԯ���H[�{������-�bH4����=*N���5���k>b�Bo/�Rn�`!w,�#��ٞ*v���>pN<l���Y@���q
��awQ��|��X�N?���Q�ld�Z���(q)��'C(�o|�ީ0L?Ȣ�Q�rZ�-�#E���O��+#�,G���Ep ������}08Zf�ك��+�ð �6}���Qo	S'�%C���V�+ڜ4X{^�wLРr�A�}���Jdq��B�Ϥ!>m�gخ���T����r�2����,����.��km�EZ2�X�?C��>T�Gt�U�����Z_4�ӫ;�T���u!U�Gip�L��C��S��S��!
,/�0
Tf���3�^C�Q�$�Ť�^��!9]�f`ay�ȳkrMX�6Q.��� �1�F�j���xߖ��0�Q�:��澀��MN2�~P��z����2Ԁ�-X�<��)��R5]b��C| #���������	æe��U��0��b�5�|��tqK�"�9S�]�¯2�D��|�^42@���GK�J�����aX|�N�-�-0��q&CwvQ��^���2@�[�l�Y��c�Ϡd�&��uS�j��(&�GQ؋p��F|�c!|��P]���-�tf�v=pN$~Zy�p���4��#>1a����P���_�*JvY���,C0���y���:�[�{RXQ��Z>���S���g���y�(���ZK�Ju��u�S�X�T�,i��n�7���7E�`s���S��؈ե�?<dZ:-��Rn
߳`q7[�������Qsf�v�
�0�r-]$�������,��g���l�.8.	��̈"gkH�Qo�5V��6���[�Y��x�6LO��/Aå��(�ߦ�F��v�n��ϲ��%>�&�_���(2����Z[���n�z�S-C��o��P�Ȋ�Ei�@ ���3@GC���4�R�D��(�ּ��pq'��Z������"�vY���JJ�Z��g+XfZ`�o��+�"����4^sӊ�b| K���o�tp��چ/ �6�I�/3
`��|zn�!͚����HW֭�7K�I��7���#���#�]�$$n(���a��>��RE=�[0m��:l #�j9�u_u��4���\5>�=�0�p�U���oMb!��!���1kaFx����ª6�^��Ξw,׳��X%̊U>|�	f���MO;}֮�_�_?�a�8���V�6)���h��Ʊ!{r:��L���=�vn BU��>I}R�S����d&��]냔C��;�&��ڣ�>E��#��PP`�o�>��	=49;ċw7R��?_���eB�5�qP����*�g[�T5>� ��!'Deu��*%.}7&�6S�?����>�򐅆W��OYQ��P�L�hm�Q�?bD��1���5�I�d���ڄX�L9���eD����|�T^�̅>f�:^,����j�b����� I��8��PD���b��`7 q���sM6� s+x"0�E�Z�܈�͗ʦtz� @�%�#���]�J�Z�Y[;R��Ͳ�ؒ��]�*�w�����(^�Z<zƿ��l~��.?��灰��5�sRk�DǛ8J����3�B?
�@�YZN�F@.%�l���o��f�[�j��9�S���Ӯ�[���\��9�'�� xB ��W?e��hH=�	8C[R!Uࠨ���l��5]��v�[�h�Oj�����ˠY��q��y��J�5` H�i�DݛR�ȹ��O��W��'S���Us��-�p�=d�s	���aH�����I�<�i�����������3���v�h��ݝ����.�
�b�c: K�b��ĝa�vob[a����	�_xЏ�Qql�����H�@�x1Լg֝��y�Ȕ����0���=bu�����-*�9��K�}�b4
on7�wY?��j�e*��A�K�w<�6ۦ���6�Pw~G|P*#ɻ�N�ƗQ7�f$G��W)��2T�V�<$��қ?�qQ�#�c�#2�y��  +�b�,O޲.]�b���-��\8G���Y+E�°�}��<U�8A�F��8��]G0�ʎ_�)�%���js��$B�nףv%քJ�Z6d`�^�ި���!ؤ�~�C�$h�,�B�Ƨ�g��f�F1���p�t����z̡�������~%�];�F�%�"���r�U�Ƌq$_
	���e������Ff.]+2X�Xӄ,w��2�n�gA%�a��T��NG�L��]�VmMf�݌x�����C�a2af��X��Q���s��mj2��?�c+>i�G�>��7u��I�#_�Y�t��[��Tf�uy��G���L�?��c!ث��!b��[/T�CF���fP�ũ10�����!���f��� Kr��!��4�P꿮����y��p؋��|?ꩩ|:������_M����4�Ҕ���,��-��ʚ������bEv�Cԛ�u�W�3�A��:��z����0Fk�b%Ks���t��<^[L�[�ݵ�s��#�����T�@ܿ_���-Jsr��7la���N0$-� ��w�T㉶eyΊy�[@�3ڱ�#c(�sdL�FF��f(~e�G��|pE��Ccy.U�Z�!�$t�n5=�l�~�b�p0����{�]aA��ʨZ���=S���ڝ*�-��P���X�pp�/�ۦ܎sH{й�$:Eb���}hJ�pi�"I�|T��L
$�Ͱ�$�A��D�o�9A0��<�~��K�V��Ky�6������B.�I�1�]�M}!~ �|c3������6؄@�y���j�!P��V���ҥ-��İ;�z@��ج}jTn��G�2|��ȸ��\�j�M�w!+�v�c,� � �uw2,����e�D�BQ�o�J���~r-m9� ��ьn���Yj̡��㌴ �1It>�#���q��o�1GOusYQ����+ϓ����3�K�4���SR�#����n�j@lѠ��[�3�MZ�Ud��h�DߖG�NG,@JV�e�|ҝ5�1��o���={�p�^�R�"����-��Z�����hʨ�W���MK��i�%KW����5���f$09���x�������#��;白�w�e�E�Nk$���|��\)�RM�>ͽwI훔�l�
�NwN3d2`F��x"��×8I�S��� TX��3�'���uH-5�93㨉u���:W�ə�]ws89㵣hu���:��G F�Fo��O�NM��}��gV,i�T��af\��}=)OU|TT��#�����%)����|��\3	�b%�=ݗ�aY	�֫
��h)�l�n4_*�l<zC�?�r�-��V��$�y�Xq��.�3.���߲Ȉ�k�Uo
��,b���}��C9�5^�^�������j�R�KFa�(¬�Gd=�����Z(���	81Nj��?�Ψ1|�,��?�x��s�R�	�ϼC��	�kH^�Q�b�ZR���Ě�i��RV�v5pL�� �ss�f�6��cm���`k�hUl��
��U��0QdgO���x�D��9�k��;�>��9�|�0=E#r��n�xX��j`�
�Gi���)���F,�E6,�
��6����&� ̃'�ytC7�`�������1�,h�bMPU�svr$ڡ�qz��r~�RZ��۲I0����v/P*U�*�>J��t'±!�2�Z�|���,Wڋ�b���p>F+�#�|P�9�o!@~��j9���� � .��E���زe���"o�@�~�V�U*�*׉5P2�!}R�B~�e��%*���7�(V6��?�v��`���mW�|'�=ݣ@��L��)m|bd?#)D�����"��jM� !o��[L����fM�@M����?�U(����^�����j�����n���j�9�q�F�����;H} �u������*1x�NE�������zT�2� ��%��V�S���+��Z�v;s����5ϒpQ��ޥ>�6��g�(?iRZ=˿�l$l�0x����MՈ������T�E�E��8kc����B�5#��`�Y��YF»Z%q(�<�o�3%�/6S�"��tG�[J\\xB����AyE �Ǻ?Ɨ�hɶ�	���[�Z��>��5�l��}5�i	vG�>hO�I�?ay���kY�uW�N�n�5��������8�����p�����X��'tXk�T��sU�?��=�{�y�aI'����	銦��Թ9��_���;x����v�~|�-����.B�㻄:���#˩�~��vp��[�^��)Uŧ�����uq�7���\Hp���pk��_O�Ӂ�)J�~���[��b64��h��*���$WG���]b�go��_n�h�w�H�K�e*��E�l��<Z��3-�>����^�w?�@|1�Oɼ��q�Qx��e� �P)4@imW�����?���Q��ȖĻ�#�Z[�}�<+m[�,�%޳['�2/��;7+��8�X�ٱΏ+����P} Z6<vnwyc;F|/�8��]��O�i)�����s��L�_��=W�$�%����`zbL��(�ԡ���|C*1r�|�Nof�(�_�G2R1��^p�����zo��wN�xz~���]�JF�
y�.Ģ��&��A���
�Qϓ&���ۮ�Fgo+S�GX�wsX���<AƔ䓧�����囐��~x0m���>�Ӡ-�z����2����e��RD�۔+,mI�2zx?�A>
��G��x�_��J��_�?��[���T���u��G�m�L�z������-L!�����T?s!�,8H�'dŊ�7��ו�!���f��(�rFU�O`��1ǁ��$��������O ��P�J�����#��2�M����u��q�����-Q�d��J���ybFъC�V�ն�Ú��1���+�^��nЎ0';qb&���X?t
���3z��і�Vjy�K,Ҵ����@��`��bJJ���v�aQhN�i1-iy���9w��{������
[��/�Rd�c�{d��e���e8(�HG
5�p��?��c:���n�"f�t���=	�~�p�ؙ�-I�<�<a"Eʩ[���-q=�]�m[7�#�V������q�R/�����i_{1x�$���E�����+��i�ʨ����i�.@�$����K�������3~�Q|�w���6.`
�P�B��#��jw�.&m~!c=cT$�<��4Q���}y��9�+��P��)E-�7�K�nH��%�����L�y��jav�(X�2}��Pҥ��Gj!9w�j#vW��$� ��2-�I��}yD_o�ь˼ɭ�	.�k���э�Q��Y����+P�5"�1�ŝ���u�'�p��Gp�tY�6���+P�ת�DB3la4լ�放��4�:�)�^��@�Ԉ�wϫ3�5Q�6Dp�i�>D �Dy�N���@�J�e6�^NR1�����%{�]����҃\��Y��RV���h�KښXAO�n�/���Kf�H�j�3�d��GqK�G��9��x.��8���3����4�^�Ȇ�#�e�iCNlĆ�خg���������U{���BnNxb3�c�`�����DA�I���^ 5��49�8F�u�3�����
���b��:�n��t�t+)���Vu�Ha:^��G�ѠF�0OT�!���a��gw�Em�(ҋ\z=�}�IlO�� T�8�$���p)6�G���F\��MC�������Bcٶ�����b)�6�n�q����Rz��!�u6r����E$$�T�n�S��w�pAp�棈�Up2�T��>_�[J�R�5��A+܉j��)Kg�o�i�����ޯE����@�eu.8�~j�������|Ew8[4����9��ʻ��$��	��Htȑ�*�R��Z���i�rV��h5Q<���Y�ߟ�BV�֗{�c��� �8kx�lh�A�vЩ0��O>�`xC:H��WkQI���`�A|���Edĥ�ϭfx��g�\
��i�ξ�*�n�gKPEw/�
c{# Y����۠��W�z$z7���:R_��m�,�S�M�-�4c�$�&�q{$�O�q���x��%�,�L��[Hʾ1zٝϔ~��T'�Q���>
=�˭VJ�n�ӱn��Ρ��Rkɘ?1���-,����)A��r��X��x%7)\�$W�����U�h�3�Z�r�ѻ���:.d��Fӭ��gr�S��{~�3k��ק�/�:f�<�0
�L�v��5�H'��=m���U��j��N���a��"}VA�:��9���&�������*O�~�a=�G��U:3�9K��I(;[�<���e���&k� ]�/c��H��-�;C��� 4��8zLz%7���Vķ9Hh'�mtq�]�9f<��\���M��{(�'U0�~ ����9��pZ�����~d�u��S��� t�_��Vֳ�7�&A��̀@2�ɋ����Y��b��4k�$�mD�V��
�rq��l�?fc�|T�v�֣t탤��	Vy�t;���h�����f��`oQ��c�	(��$��Ձ��a2}t�T�����#�����BG������
�R�� �}?xvB2�=O֩�N�*W X�X^`
���o1��̻�g�dW~H�&�`W�\���E�+�`1�:R���d>	I^k��M���ڼ��^.{�1�qvf���rZ"��C�ƾ�����3
����G>f�-��:�w�[��])��y��Y�&y,���=��D���	<�r���S����.���L���N�����L.�@�T'r�d=��Z�p��#�>��Bc���ӿ9O{�t��i(VP�	��Vn�Z��̰Μq�/^�a�=)q�&�����;�}���3�dk�����Us���tȍ�&�i�ؙ8U�Wb�t���!��<sX��i���8��%M�Ӝ�{�?��_���Ujl�q�|ڛ����MJ=4�C����K�'��3��
��s�&?���f ���4&�UϬ 'ӽa,;Ցy������\d���Ƥ�4������ �X���צ������s8�F֣B��D]R��{�`���^��S�s�)�2�ӿ샺�'቟|۩�	`��2-P=T컻Q�tY_���R������2z��J�xOB�d�#�[J��E�z�a�|��sj��F�+B����z�T+Z���s���K�я��2�q����� bYi�!Q*�}�/�`A&�j.J~������nW4<Oi�9b��ѡ;Z5���^C:|De`��&���o��.'�1zP���ӒqCkd���N��PT�%�_^�zHP�K�u�'��LBPAO`Ϊr�p������G��e��w����0x�4M�Bs���0W�[���m�%8�1�U��g)Isp�BS ��� ��x% ��������u�p^N������ѭ$�k�)+N"�d���#����^j�bC�M�p=+ۏQg���wYYx̐����05���6_�|붅O�j�"ø��O�.S8Jf���������*gh��àJ���WZ�V�qk_�կ���|;w�[�$����І�l$����J_?R�d.���V��B9,����}ln��?�s�|`�݂D:��X'5��9��~]/i�׊�gF=���p#� ���`U�j���+�1 �o@���V>r[��e��$����dc.�,% �@�E+����SL�,z	��[>��x���闿D[�К9�#CHܮz��߳�j���+cs����`#�ǘ̴6�3�XS}:��M`bjr�5#�y��Gf��
E�7�.U\{��C6�hbs�u�^�{fV�|��.A��j��@��_v�n�}")*n{O�^ B�3��o���U�N�����##���yr/���C��{ $U����@'z�#&%/)���S�\�G������f�ew�<S�:]�1�/b�E4����m������	7:����\<m$����oE���[� k���'�	ΝuN��!�7mZ��a��!u�޾!���{j�����0t��� ���A��Şh��o5Y�1��۽��%������mt��R����,J`��+L������E)/�Qxڎ�V��VZ`tJ����l\�)���2���:�I����s��D���l($U�q�a2Uy��hI��c6�V�����[_~�qcn��ԗ�CǸ���K	��Lͺ���?��5� �/[�X���i��K¹��OɝDW�\>Z%E�rf�g�Xr�k}�C��+�I���3�����R%8���?T����*L�����s��cj���۵�c�EwB#6-f��Dl��Q�QD��42���*�܆,׍��A�"v*}��f���v���hH������)+*7��=���JfK�K���x��ݗ�A��Ia>���#_�8��R��l�~���N*��A��|�tRu�б��cw��<L��J$R��_P-^� CgI_}�X�1�Ǒu�,���P�t�w#��Кg^f l.�%�W������A�WxZ��t��+%\�$��
�i΢�w/�8}A��O���A6`<�^;>l����]�.ID�����sE���i(;jxɂ��U{��q�mk�r,?B�_�Y6A��(��}M�p*�.�>l��*��c]���"������w6���n��[ P'64�*r��}����3��D��Q����������-!�>�`�����xjx�ܪ	B�n��]M���6�t����Ø��;�{���*S����h�X�6�[�C�H��Dgz-W�17�{�6>
b�զɱ���`]VQ��u��0�>�E$"X�5��f�M���W�j��BP=?+�� ��e�:[5��=�ai�r���Dl�~:Ɇ��6YL:�NV��}Ld���0��#�����gv�N�;�{tz]�>a;
�"������Z9�0�&�r�K���2-O���a�����j3��o�6��;H�4<2���&���U� �:�phH����z��;��y����Z�LG�:l\bV�F�H��m����J{9�S��[���2�O�e�4��+����&�Rp��������ϴ��S��K��*�G��C`����9A��8����X����n���t���
�2$m�H V���?c��OB0L�0�)9�2�a��x:�V� ;trWhW������6��Q�E��z�(J6"��%/����}�Ӗ��y�����p+B4�_�"��
�����m}��SB?��O���NS*DW�����V�
��1o�^_(e��޳d��s�W�\���r��-�{1&����"id��	�����"��wM龭"�H�1e��v�r9����/�@�/�ξ)�ѣd���Tmb�T�%.���ӟ�dՐ�o]V)����Ɣ�&��dR�=�������	�eZrA}S��-�y��t*�J2?�P��9w�@T�Rr���צ�����z#�#K̳ȅ�<G�&5Z�7��=�P��ÙÂZ8k�]��q[�^���=�Q0&�����.��6�@Lk��t�+&�s��tU�O&�pōz8�l�Wo�U��-�!(=�sEY���ޫ�1���> M?���΀��ɥ&;�WƬq�e���?��ƕ�M�����]�4�,�;'�䄨2�)ڠ<�?�-�����`�4ӟU��'�Q},��y)�⸾�ѝ;�Ӵ�4e����
�E/�d���4�\�+���F�p�ӧ��R�*�M�`�몁���s��*���J���l���/ۖ�R`u��-}��ۜ��r��+��r"���rz����U^B��#g��d|uz�e�)L��������b3B�)˧G�(T���5R�b�n���V��_��e9�,L, /�+iN�v*�8Q��ϣAs(.7]���B�tWP�iE���e;�̺T��C'�OD�YW�Sn��V(�W�'�)�P���� �oCX}��c���8X2T�3��/^�/2P���u�S�9��A��u��u�w���̹�ȹ��@)�������x?�A�G�@�⼝X[�@Gb~%����B���TXI�)����; ���d��nr�G����S�u�s^{#����i�`�x�7����"�*�pMQ�hX�^��C��Mp��͏^��k�CY�鿫���0�'��cF?�I睅��0�/+X�A��{m�JSC��"����Z�����VJuW�;@V9��_��D�m�Clw�Q�$����#vl�����1_,�d�R����_�_��9������5lC���i�����F�^'�;9`��~j+e�Њ=v^*dOFx�J�����5�ר��8�� ������
+琘�)�e��1$R���ц�.� Q�Ex����/����z6![�o�����7��S,��,�ʖHixz��߀�Ɍ�J�+p~�԰r���%~ǅRn�A 1�.X �r�fȤb2F���7y@�-f�԰E~>A.�4?��!.������s�͓��Z�{S��|��h.n��7�:@ug`_�*�*�)^#�{<� �*��
�/����UW ͖$�y��֭�ڎ�]0y���)���Hu�Uz�>ȡ	''&r��/�n���d�G�R��M�ۓr��< % ]�!-/O��48�����U�P�	�b��.<�d��\��\_Ö-q���	;�eN�����5Z��c��U��kpG��`{7�w��_<�=$>�1�ؑRu�㽖�h}�@5�a ��f��Lc���)z����n>�?m���J�B)+�Y�W�ÂRS-��㝎68ЗCe��jbJ�4ۯ�,:\�E��x��|QŖq���㜞�>��C�(�qQ��2b���@�I���6~�|�߅�H�_K�q�aC����Ct;m�b~�K�p�L�������U� 1x/h%�X��N��j6K�8/Л��qE�\�h%��Wf�B^XR}����I��+�`ot�Y�
%�:��L�,�E���j��M/��J!��v��0�Hcǚh�R-����1�uepQq:C�] �n#�,�N�*X���U�i�}i_[f�r��C*T�������sڰ*O�A�o�W�H�YfxX�K���x�{�������a������8*k`��3�Ӥ(��e�[s���U���pRb�y��%�٭�	kq�bC�R�_��2^�g6������]B�	,� �@t���?�4gKj�l���N����A���g&Mt`jr����~���w|/��AK������>7���Y	_�2�[�������J����;(襉�Ͽ��0ʠ(�m��,����dF6N[(.<�M��$��{��W!�c*�(��Ei��T��$��#�r��p�P��ςWv��J�����3�"aܝ�[�;���Գ�q��! ]`r�v���+jf��W���V�1n��4M6�I6;�[��N٩0�.�H��{���w�M�����}D6����D�H�|g�����l�1�_1�#ǈ����A���P?]���������gX���]"E�ہO���z��˺�]-�"�c-/��.��7�쾸���b<mO�%��x�j�Dґe�r�7�>�<�uN��N����g���+M2D�i�����c��DȞ����I����VK�k�ئb����{����wA�rꛃɕ�Uu
�q���樃��"���Ppu&g=��_�ŧ�����x������7���R�q3�G��:�G���6��Sؖ��X�j�B ���Rޏ�����d~$P��ʬ��̈́�2�7���.o��^{�0��]yDV�:�{^��iYQo�~>�M$��#bug�` yK�W��NMK�L��`��S�MJTBa�� T�ir�� 7�z�`���=� S�Ga�ã���B�dUj�-=��nş�`�b�^���G�QL-�i��+�{-�d$��X��:��� Sc\٣��a'��?���k��lr5�'���5zY2E���a��o���t�>2��wr�v������n��ϭ2W��h&�L�� q2}��^QռڇnI��Szzy� �n����ȥ�iA�:��r�@� �&Wi�M
�B@"�w�rȋ����DZa����"�f*�����Z[~Gg"p�f�H!o�� �M:"%_��̠�4��G�E̹|;{ɝ�?oZ�Tt���uL� ���IOȵ
/w|���!H��h��R~�H�7F`�I&����A�����	OC#xV�$_���\E��M3�3c�}?0-^ѵ��#���<�u!�\4��q��N�>��X0�L�UdI�J��!	�Ίha�k\���a�e��y~��"=׎��XLZ��������D;81R�z~n��F�yGܑ�.))1�h�*б|��r��(��r�\~�vIp�U�M�>�/�N�P�;*����*���J��2���>�%#��P�P,o{:,�$��9�ȋ���O��݌����me����,�6��3=�0�*��#��������be���*�?�7Ab�6�~!?�~'����+�AW��v�����CL*ǗmV	�?=��D�o��L���D�/  �?�LT����F��ZI��I��MH�}}^�%�.�jr������;����K����ו�K ������P���x]ӴEhe��7���
/Cp * �%m� �m���KZϔ;M7�F���x��������(���Z�Z����lّ�m�1�I�;�b�§��M����8EC�'�!B�sd�[jY��Fܓ,%��4k��o�M���z�Ɖ.}S&��N��[d��\��7I6��� ���? J hc��	���[-���ۍ���ogl�:�5��v�f'h�?�L.����Y�~�²���515�j��$� *��B���L��J����'NZ��n�.s��}٨=� O�^�-a�O��� ��]?�$o3����9�^�����vV���)���c.�AԻ}�":����=�=��}v
��[\�C ����Ъ�^q��;��l�H�g(o��ԷI��ރ�>��F�5	bPV����7*V��z���QFb��o7N�n���w4A?���/*~�S�F=�<tT�aoK�؁����wYʶ|�r��V�\�	pQ�bG�<����)5/�&�ww|ޱ��?�Q��l�#M�W��+�e�,Os{�MT�;�� Å���8b	ً73+ �Ű(r}�Lx<P���d�F�SY8�E�]�Y��i�a)	��i�s~��fr��)�׾������5:�`��4�y���[v���C��|�G �(�x�B´�gE1:��p�>���z�� ��K�R��~ \�]v�bF}厧�s�6�j��}��3���lc���S`/��sx��?��)�Y݃8k\Q��`�1�ڬ�\���O�"Gb�Y�R�R��+w㪭+�3�ǣ4G%�F���&�^�[�A�@�7��i�Z3�׸���]�D���v��N%%@}?�e(��Ґ71�)�r�?{�Eѽ���b�����l����hd���
ќ�`O/��a�K�qA��E���y~F칪9S(�x e�j܂��f�n�e�P���B�eoNx������9iu���q�X
�曇���]��N*]�3w_�`�t�K�Ш��I�k-��X ������Ȭ*[u��������T�:JRB��o&�&�Ȗu��_:�#UG3ĿF.O�%��23���gi����w����\,�S}�d�Oo�Tp���`.�Pp)hxP�O�g\f��5m|�0:�ʹTM������)�n���Ps�zֱu���L�}��7BȆ�I�ž�����b�Dҕ
��UU"v��v�poZ�l5�i�s�NqnjI�KYGsݛ��:��ʣb���,��H�8q��j�=U��P�|w�e�֍ī��	���n��;	��dHq�y��X�Rj���T=i�K�V�5�"ex;�Ბt�:�	c�)�2�k���l�L7A_Lh��0�W�O�$�x����\�k�db��Q��ͶW|�d�E�('�A�x�ӝ�e.
L�i�`��
K�YôE��x
շ���{���"�݆�,��7�ZE�lڶ�o�,���M� �f�K$-��q-�԰A����R&���,�;E�M�c�L�A^^��L �?�9��>|o3�_�gJ�����d�@�	�t�lk� �q�߷
�S������ӤdLXBV�%�D��s���+�m�m+���z�Ork�J��:��ʪ��&{�r�<	I�~�@M�
��>AD:���"@�L�j:끙���/Lm�?IB�3΃� ����a �"�"N���=9�R�&%�e0�k.O�Xqao�Ǧ^t�3�&2����;��\<������- � ���H���[�;66�� Z��t�7Ll��170V6z?H8Zmf��ڏ˒9�b�Svz�����0ڙiB�0�U����k��p̄�s���$���~SN���4��* ��0��MIAD)9�2&�ɽ/�Y���)~�&�;�VFym��V���d�J����pƛ.�Zh'&��:��]��V+�9;�1ph�<��C�;K�Q��7y�(/���oɞ����}�l}�X^3������By���
7ؾ��;�}q2B�ݳO���N��"W=�L��G�
?��o#���һ���d	3�]�WBw�\��}��t��R��1���3�d�p	;������\h��2�m=�1*b,vs�>���d�0�q몾��3������﹆�3���xg���)���[]��������#&빩in=�����Ы	���r���S�%-�>T��9��O�m�����~�@9*.rz���T�E#Y}]̸N��U�kP1��S>�P��.����Z~&��bm�q�v�^	uJ=��&>d�H���+ޥϟk��_���s)t:Y�&����He8���W��ۀ�R0!�Cs����ۡ�Ŷ���N�M�S���,��A֥�Ֆ��7q�=��M���LM|�	
���'0I��J�%��?�����
��+8�4�c�U�;�'+�,��y�$A�����#�8!�4j��ٳ	>ƊfťI莹���͏�� �FHruӬ��R��ے������(/s���dcc�^�E�qVЉ�����*`Z�\-u���#��Ew�_Wh�w��xfnz�[�ꪢB�.�#�[��)DSzc&��.��eX�Q�0f�MBA�2�lv�T]j~�m���g�Ƚ=(��A���n�� T��iD�*c#^��NA@.|i�hm���@�W&�Li
n�Z��;>,���)Cly:D�����������'Y>1P�//�ŃC�s��HD ����T�?C�`�^BٵP�x�u��#�~cgA��ɪ$�ԋ��uGR^�-� �E$�i�@���&x$�	��	oe�H�b�"[ �g�+%*���dT��R�I%�Ɉ4�x� pk������F����Yu���^ ���O����Nݽ�۟�"�o���ˬM�E^!C��9po�/��_��p~�Yj���M�0�d>��Ѽn�j��E�ƔR��F�� �J�l���8{\�?�ԙ�Jh1�Ẅ́�V��%_�t��Rnȯjw��$���Bul�C7��(_qWd��/������^9^����l �N1&��#���m	��R''	�9%��~Ϧy�t��^oaA4�u���^�ˀ4؜�����X ��C�~��pY�u��e���$w��햓_.WcZ VE�EM�!C��z��k[��Ѻ]�r��ځ��3�U&jH�M�z3��ߥFU��A�+�M�Ե.��Rb0��#h�&�d\e�XE匡+��b�������y���f�vEcM�. o��}[�ڮ��1��s��'�~A�{���|��U.�O>\� @:=�_�و/��)��{�6� �c�͏ ���}U����6�Փ7��k"6y�:l⮽��m�	U?Uo-ZR',�c&`R/7�t���$�G�X����=e<�]�\O/�ef4u+�?`�u��	is�l��<;��	��Ρ�,�A�6������MF	 �;N���%�Z��(�1��Pؖ��{\���G�Ǣ0g�6k#��.����hb�35�i��j����+��ħ,f����п�z�/J��+>J��	������;�ۛ.��=�~K�JZ2��ڻ\�U��I��Ĵ��;�ϗ�h����R�w(��q^U2�}	�ƭdI���6�]����b�_p�q��I�F�yCy�}�a�K;�qL�������7ł�/ͯX��O�["RK���Ѐ�����\0�1%w6Af>bpX$!�}����]�I��X���J�~�%jv걠�Jݠ�[2�I�S�l�زN�m;�Noc,���-X��v�dZ��Q�*��&^�3IU��������~�T�"}N��fY��h��ٚp��h�x�M*��z��¬�-vMf��'K�ox����g�q��ɂa0Y�U��8�R�����Lj�����`�n�lR��ұ�X�)���.�7�'=[R?�_I�^�=�g{f���1A�g\Q,�C�~�t�PL���g�3�l�!�	}���lA�m�̂teS3\��cc������{G�J\h�^�C�"�� ��?�h
��	:m[�e9�"u^��?�l��5�(�vh��h�=���L��Y3��ىi��!�5��2��(��lڴ
B&�.���]�'U]��U.�sv�����=fO�G�Q,y�a
�U��:�鋸��&!z{q��G��4f��0v}MA�Zs�
.c�D�$�:"<�ä���v1�[cV��*IH��B��QŅqn�F�U�KHY���OԾ�������Jjп^�����b�1v�	=�*}��؝��"b��ko�ڱncw�����c�*�X͏M�p<[:P�(Z̈́�N�R�/w��U|�h �}�����Qy�j��Äa�i)����=�����؂�?�:5Q���#���ޚ�+�a,���t�[�����Lg�8	w_��V+��X�o�j}���<W�zn�F��\8_e]In���]T)P�U����s��%Ms��9I�e�6ֆ?�ߜV^`�1�����rB���VCK��������ߩU���g^1a��p�˘��o�z�Ǟ�0��٤~gf�]��F�%��7������32�
M���`�|kF(M�+4O�X\�w&�j�0>�A'a��(��>�v�\�_�4m�_��_�0�n�q�E|�2Z+~�k����u�cmJ72�} ?]W�>k7G+�ȹ�����_����ݙ
T��3u{һG�aLo���
�ح5-!���
��T�{���H<樀��+jq���t��!�<Af:4a���Mr����mT�҄�K�f�ļ1��{/�pƔȺ��p��9��|�MhW���ZU���S-�]��S:��,YOb�C֢-շt��h��ĥ��2r�ﰎ0�+mb�>����t����O�Oݷ�	���f�e?x��@ފV���J�ȼ�;�a�tNZ,�-
���3w�n���Y�o�[w\ڳ+acj�\d�2��������(�ԬG+A�pό;���c�n��*����.rt��-=
��~4�p�������*�a�VJ�jUk��_�=���@���)A�1�A�8�F�Q�2�/���H}{R7�$�G�Ed�*$���i�a��~k��s�O��$_y�F���{	͕X�~��;�X���6OA�Ñ�fB0���s�W�ϯX~� �c5�֐=p�U���FT�y:Hˬ�zPI���3���D�o��F��<�R���j������2>��g�����j:��w�9v���Q� 5�>2�D���D�@�49ӌ����)�����~��Nym�w�Y���ⱌv�1K�E������1w�GQ�Y�{K�K�+���ز3��4v�l�U�+�J��*�g���@.�'��3&3&��D�*�D�zE¤N�gE@�e�6���/�1@ ���.{�[�EҤV�ߚQG�\Y��3�hh�n����Oo��HK�2����S<���4$��*�9b��xO�9W:�T����|l��y��IeE��N-�&�����$,�� �y�x�� `���lN9!+3f��`�xB�]��C�I��߫g քU��E̬��u�"���Ј�K_��å�:����&��5�'��"uͨ�:�G�5�Fq�O�6��an;���gXEc���I�J\�Ry}	�OR_XT��\�堷���!)7�)��[q\�R����	���ʶ����`()��_n��U��A�zER�0��DK��=ߛ&L��U�n�t��M���q.!#(�D�$U1������?�����+�5`���:�}g]jX}�KH���j�4�ɯ��YϽ�����u8�m0j��i���|F��|��:!��u��K�ļőV	���H`�B��uR��\�Ci��Va��5�LJtjڜ��C�sָ��c/����2k��bl	?�P�NW�0��O_�x��T���k�+��"ֽ܍\|�dEe����H�x�z�l��
\�tiC��뀁�H��Ex�$
���a���^�hb��N��;%7���;og�+�,*�MR����$\��q<>��0����Fʺ�s,4_�Ѽ�Y�� T�pN���������>+�����J.���2f�o)/���?k��1�@�7�����+{���=#��e�Xq�{%�ձ�bib�����2�E�$�'�reKJ�y�	:�A��A���r���آY~N��YBTm��:'����[L�9��0B���������瀌b6��)#q�a�3�"�
��{ճ9��&&tF�_�g�z;;O��a>v7��3#��J[2;��S<F���&�9�Eb ^q�lHC#���x;�q��/�獃�L[P� �eV�H�rm�$�����9 vQ�b`V���*�s��HM��&�"�_��&p��	��j�K��v�5S�pi�X�m[�+������/�ASQm�!P�Ɍz�)��2����DF����m���V���SvJ���`T��c�ׯ����J��L�V:U�;�Y�h�6������ �Q�Y���(^��~�7��r�}u�k�}��m�1�B�a�6o�
F|���a�}@�BS;�O��Ng#?W������8
N��o�*w��V�d�Q��eW��M\���W��A!1����n8dZ�q	�j��F�Ջ��A�\�1�bBv"��)1��7�X)C�\��� �x�5��.��h��E�����|��x ]���p#�Z�g&�Re�;=���!_@	��r�5�S�EJ�r������P�A�͊�@hAr���׺��q�r#�:�G;c�#ӿ��^��**�BP���W�hZ-|���xq.��^X�j=�4&M�������~��Td�kL��?�sx!�ti�Z&����dN8V&�W��{�)��!<~&sټ!�
�Q��|N���M�L玜?ـG�,�:P��}�q���\,h��vMK'd�m�K�@��'�Z�F]��4}?Ӏ ������D4g
�U0�='T�,�8y�z��Ҧ�e�k����4��2�"�{��˱�xa�ȰZ�&�tu	F��0�;�RbU�������َ�9s��i�37c��?� Z� ���*N�`�p-�h�~�ux9��p�ݸ���z$^.��oB� E#{o����z򙇽Z��Ԇߏ�����BPb��[	kT,[���S��^����0�]go��T��ذ C�Ai�P*mk�p�A���.�
������WC|i�0�	,;��t�hD�C��$DL���C������'�PH��4��C����wK����*T�����l^��P6UuY��͟�A�m��3R����
���=1�����x�1�lxSS��4�T-ȼ1��[Ϙ��ؒ%�T���^����pI4�I�#���������X��[%�,��u%�f^����zѮ���/�j��"%�"�ET�|B�^+	�C���p>%�r�����Y�����0��X���;�]z*�P�O�C�U�ղ;ݏj�J�⽩6�G���G酣�=J��W\:�VMZ+_3�l��mהw���$�J
��s�le΍���_�7�dό��M��s��9-y:����l����|���6��#�$��u�'��9���~~#^���Q�u�Sc(��ޫ������kB�Ld
 '-�����*���?e��$f!��etq.^� ��E��ʲp���5z��[�c�����ƿSJb�1i!Ǥ�$H ��zB"hߔ�d����+�Ƶ�D�D��������U2�k��X4�I���\b1N��v��yTW�f?h�E�D�.�,���ԡ����ݙsY���퟉{�Ó|��.��K�E@	��_��U����)r</{�AB �؂͞���c�U� �8 )�d�x��Ǆj��yo��w��\�Uϗ��'��&��E/�RӰ. F�}1G�}Y��_O��0�<�g�]��b/��4L'�.7*�d��	8D��(<����xUI��*:�p]���1w���e	�JN����x��Z�)�5!�BP��	�{K����v�Q����ܑf�f�Q�bh�q�5���ᗽ�@j�ڹ��Sl=�S����cJ!��+-@S���f�����S�J�B��@w��gJiE���O�\�h���QޤS�~Ū�]�KI��k�a��(�]q���2v)��UϗI�6���l�ܳ�__��qd�Y��؃C��v��K�H�L�����������\/|�hX=/Z��s�KCd�ЯI'���\;!%F�f���X��$}!��}�I����#�m�>%9dJ�`H���z>�~���� π����$Y��t�ܚ�c���L�-�9����3��Q���L���@��m���<���}}M�fh#��W�s�i�Y���h*c*���p�\��f]KK�[�x��`�z��$�za��߳���8>�aOt��t�3��o�Z������ExR�'G�&��8�������d�R�`_���^#�2gʑY��'�P�DV��,����-;t"���S�g߉�l�"-������A�S{"�t��u�d+�^�d��c Z/���A�8��ʱw��w��/s�2�ﲯ��m���Q2� b�(|��㸶vL��<8�m,f,  ��`*�6b��(¶�M
샺����/���c>�B�#_ʺ��Ǹۨ�7':�k4UP���n��^����3�B*�1�H�O
j�h��ԅ��!�l�`��$����j%ZO��f�j0!ndMJ�/6�J�����ī��\�{V����/�F���/�6C�2��H�g?g�1��C��1�P���������g�y�ȫ ]K��
��qڊ����"�`u�cP���W��AP]��"��/P�.�*E7}������,�O�(J�jU�"�xD��^e��D7bN<�w����#����<]�?9DS���?���]�X񢞪B������V_h+㥚^b�ç�cv��!K��ڃ�.��ֶυ��z�Ι���h��p��3=\n�ಯ�;5|�9�����R�r/o�)��R�]�3�n��ο����W���1����Z ���Rrxu���d�Ř嬠�n͘(R�˲¤Bi��0��y�:�_B�*йQ�2�>I�8צ���g��y�헾��Ke�t�+SI�zTV�:�n�}�C�?�7��`"	\Q��S�K����.{Mdi�r-ш�n���` r�/k�{��Q`c}�����?-Lf�Ԍx��MP��������ں]�Uz�w�ak�& (o5�\��I
$Y�yk���P�%�7��m1r�����֦
�q��{$n���������&�����82��Ż��S�,t�n�puS����A_��L��9=iUl�n�@�����=�aSd����֋�i�&��GrZ�P��D!"� �%�9�Zo��g��f��doQ-��a4b"�7ԇ��S4M.��Y�f|�}����o��t��x�	y^ �n�I�i�
/�|)�!\B�<�+�#��:�7Z��I��)��\4Q��L@#�$s'��5����A}����0�\��Q#ҨĢ
u�!%4�,?�K��>��`0���Ux�r���!4����kp������y��%�-�'�"'�X`h�����윒J;L) �y���Rקh�ܥڂ)�U�h�ᤱAr	��P8+�p��vݳ�U��>x���b���s��n΃Cnb&�����)�x>t��#��<P?��o��(���9�ڱ���c�%� 骜��}e1<�@ �n~O�D�7*8�����On��0��ed��*�[;7� m6��?d��λ��W���H �����L���mjN�?ђID�It����X����u�SD4L�E���_���۽0������пUc�^�*��°�j����t��OcB�gD��_.��� 'ש
�  �x����o��xq)*E�}5�[͆u�C�
 �b�%�K�.t��oZ<>;a͡����/��R�h����(��>ZkD���lmǂ��Q���X�v8}�j�O���?�s'8Y�݁�[qB0���vY�#DFpǎ%߉���do��
�JX�Ɲ�rS����b�[�5�\�Q����/f ���?4�^h��
	�Vf[��\����G��l�]�5L8�v��Bh}���-���:%�Y �S�F督-c5OD��8+u�����m7=���@�;'b%���Ys��m��=�U�t���V�aw\i�ɿ
�8�8�8#]g-�M�Ůa=��[Vv���� 鯖?.��*�&J:����xr����v�d3[pU���)i�.9�>�aq���Â@Hޭ�����d���$�ޗ�Ь�8�I�Hb�} ���*�>j�l#Ab�]o���n�B�wȼ�����*��Z [<2��uG�l\���F0w�d|�4�������Q&ܺӽ�N�!)"6X� %��?�E��?���Q����2�#�x�k�+�,c�,�� �� zl����Kt8���ٟ�X+�k��<?�}.M4<d�3'ڂF�{�8Lp�]������)�Y��Ues�r�;R�=��RF���y�ɭ�`��*�����~�}C��_���(<�O�։p�!z1�~�p�,����zݟl�,�fĦ~�wE]�>jF6��U���o��$�S� ��
��^��
�I�RF�z�+A*}X�ws�q�ZxA����U�60��WԤl%�m<�O��}W�[�r��R�2�Ӑ��!��Yۂ�mm�-V2�I?J�c>�*OG;�
Ȇi�x�_��cB��*cxT��Zu#�G0�L<�(�!�غR!Q�h�Wi�Tm����տ\���j�L���z�!�J�f������r4�&������&n��q^��%�_�߽�~��%�8x��f�؀I �M�O��z��!�߶ �	c-?�������nbt�#C�e��d�;�#����Q�L���di0�D�bTN���u�t�X)-Dʼ
���DN���$�2���J@�����1JB�w��y�a?�N���-מ����w��X����Y [�Q$�@d$c��df�qL���Ѭ~(mmGx��p�r-��c�E����P��t�S�=��]~��$p�.�e�.�a��u�����=B��C���;!-ni����ʟ�f/��<�}��{��w$ʖIE�̄3�I��~i_��7�;�2�$L�k��䶨�*�%�~�l�ex�:��6���~IB�>�ˠ< ̜-~OXAcB�d���¯�_��3z�y�L��F�P\<���%dy�|�O�)���g;kj�Θɖ{(2��٥�\%j�K�w��vEK/`� ��2[���B�D��5��c�����?,ܗ߄o��ѻ$���IYY�Qgr��c6-1�_�:���|d�?�G^�Y@��Nؒ+~����3��4C��h�"�q�קs=w^@��e�|3;�8��-F���D���}N�'@�HQe$�r���1f9��M<{�h�M����ڝ߇_��$��`�{h`Q���V�\�-�XT�KԳ0��T�D���N쵊�9�x�T��ł�����t�L��;σe�sN�����%���q���������Y�N���3s� `5��G�Ĩr�5I����]� �[��b�Q�&�u7���F��8~`�P�h:�C��?�dY��U�uz��:̑G��F���O���.?�"�ge}knP���2A\��=}�}�O��Tl�c�R����3)�z�K��\�H�1º�.�Ͱ�t����)���n������z�BG]���ƶ�~Û3�+�Hi��:��^�%N���U�������Y"k�u��_5�rW���J� j���KUns�����F9î�6��-}8m,+j-1��ݳ:|�UW���'(�����xA5����	F�UHmC��Q�^)z|t�:� r+3qZs���T͘���� P��%S�V�E���MZ�_�;3�OͳNq�0�����ɞؖ}�'�(���Z��L��-�l	�^�o���H��|�j�F��/�8+�d�͏�B`�Ѵ�):Y��wF��4%1A�e:o�t��\~����SD���4��[
�\8]��zz ���?��h��	�M9[�w��A�U����lum5^B�v�;h����u�L��YR���ض����L5a@����FrsT/��.9dW�tW$P����H���g܋���-C1?��X�l!��HuZ���]7rӞJ��M��'e�"z0́$�������!]⪌"1d/�-.=�D7����	�׹�O�Q��=���c�,D�e=��7@)<m�I�pqC��s'�ҀWwD����?�=֘`µH���q����Y;s�V�7l�R�bIgY�v\착��V��ސ�
����@��G�=��	HpJ]D=�,�����\���j\��<48��e"����R�V3��.���3������<m�1����Ե v�xRS뼷��Rd31o,ˬ����l
G�� ��{�0��"y�GR:�����CQ��>�g�#�׼yg���y ����KƤ���|S�v�T�kK�~���V7!��`�w���#S+��ؘ���2�djH\-�{�nW3`��Ʌ�>��;�Q!s���G�@P-m�|���/^+����1����к>J�̘�k��a	�5f��FV(
|+Y�#a��l��F2?��-�O�8�����1���n�x��$��54&�r��<{2�X���D��G�n��S�����		���Ț\yi�L���^�@W���$_�b����>���z�ȀKL��Z�RW��y�"��|!U �ZpVZ��g~fj��o�?^�"�."�v-���4n�/Ӛ��|0EƝ"H�o�ët����u ���Iv�
p�|�xV!�������3ֽ�7[�0I�rz�G+�������#�;�$4\��K	�#+�b�U&�0"�t�J�#�X6����u���4���l��>�uy0��U�eA�K4!ޏ3�ݱ{kqJ���oºcI�n<ή2�ßHX!�d�e/�z	����;�.Q�o&MOQ��H�o�f�f)���h�o�1�'rJv&䱶 ���/v~N�U���>Yo�c������	�ۃ���F*�6@I��y>U��#  P`&ko��E���9/v�/db$G��RV��f�eRa9���m��oV���*��{�dUj�0(��1��e�h5*5��76��6c��?����n��W��iG����LMLm�M�?r��D�-<����YX�ω�ڔ �LI�I�uPwޏ�'����d�%��v̒^<���#�Aj��/�Z����HBT�`�Ը�8��H� �����y��!Ex2��E����<�ͧ 	�r1 :�%�꒢a�ZjZ�۱;b����ؒ�ӟm���	���(n�eZLF����l�t���ȴ>Y����������TiT8ZhW�ܙBO2v�P�gYj�^F.�%����~�oķ��k'���q�S�R��*#[��^\��<����0|� �(k?uFhX��	HϷ[b/��x{�(��l�.=5m)�v���hީ荮B��۾�Y�n��'m��o�5p�E�y��G��y�珐�?��g�h'c�v�#sD���M=t�G���aX�k���Q�Y�d�yK��1�������bv�z��1�����.��r'F:0��rVtĭ�v.#[q[����r�o�FПW�q|���#/�H�p䪻��ۦ��{X��Lp�_��ʝIb�}C��)*�{R��-bD��o,Ihn C�wiͥ�z�g*�=��[YN<)��۶�J�͡}�`8:w���|`�<�����j�QG�2���)�xdSA�L���&D�?�%;Q�Y˖s�.#B�Ң�\�+� z,$���°��!&S�~���8W�K� ��+U���'�}N�<e�H��F+�p8���]W��ʞ=g)��Ēާ3s� ����~*�׳�֔���j$`�p��Z���A���)C�\��<��B��w@�v�:1�rTp��X��bBz�����L?~5�]K�FF�z��6R��p��e�J��~n
#��u��
��Fv�+B|X�*{w�[V�~��A5e�����> �>Τm�m]_��K����S��2(�Α�X�a��ۃ4m��2)�7?���>yw!G܌&�G� �Y�<_�����ūkL�T Lu�`�G��L�_���ػ�!r���oT��z����v��Źa%�-����!���f�BB�0�Pr��������`*����\�����������	ѩ����w�
URM�c�<�⪣ d!<_y-����!B��Z�bU�7C�?;Յ�ΚC�����ͦ���N0V�+b5�����"t�AnS׼k���1����n��qC��w@�良'�J�z��Bwa��WN(�-���ٰ�w�(��ƻ�Κ��[P�o��)�c8�d'��-� ��J6(���G��pom��#c���
a�1�Ht�b�=��~�p+jՕ�{�ƢaQlqʸu��!=c�n��:��Y��z�԰�ʀB�/��Fܞ	�{��$+t�ErV1ԛ�Zssi����x�\�ò�B$����T~��IoT��,X~��3�fK��[//6�w�ߙ�B>�K�A��]}�~0��cC������8ؔ�#yz��z3�P��~!%�&?�=d���H؊����jď�W-�2����, ��B1j��Qw1�Vv�O��ng å]2<�=����D�8���'��ZFJ��n�}�4�0�ќ�
���Yz��~�����1Y��۱e������G_	�Ya�X���f+�m��*�b3��4~�棵��#������~�7@|�
��j3���eԾ�x�_D�J��eNW(@ZPUe���ҭ�1�=ɚ��{�4�n@E�2����7a�j	��]�h!ZI�g��]��y1�K5�������Ԕ�v�'9�y�x�+�.r��K��K?��ͅ���ee��N{�ï�G���R����N��3�������N���3t6M`V+��ju����I+y��� d(��C[�'�_uX�(�I�I��k���;l:gܹ��=k������u�7�:��G��F��O�|B��m��gf`���R���\	;L}��O ��T-TQ�3 B���)c�� �\C���.��M+��qi"��E��)�B�nD�l�-�zS����r�Mն�x��4���#>���3�݄���(� r�қ�U<HР���O�_TI�5n�}��&�ʹj��$KV���8�ۢW,M��ݸ�gJ��mm8.�#j���<�|��
�^Ĉ�僫�����SS�	'��Hn=֑rtR���Ī��i�V/��5����r��'#����F{c}
��.�k�&Hl�\U�f,e��0a��O��ux�N��k�����C�*˃|�sE3ȩ�~+�xh|�z��
*r�iы��9,��V�EF�{
8��`s�JU6�Ԡ�3w҉&�7�T��	7��i�,x�RM`ѳ�tY$�a�q��R�>K!�O� �1`D,������o��j3������砓���~�>����<��J<�� >���Zц�1(k�&�ƷG���yՐ������[X�`�%F�7�pd�������p��ݭ��ar3_g��:=�����5�r<K�&�~\�F�'D��%�:u\�HLork뾔O��R��
+�\׷����]D���a�Z>",���~9�=T&B$��\����Oɺ#a�Ʀ�I�3l�_�X��;���<��{�tz$�&� ,��NH��霠�;S+�����p�Li_N�r�Vs)H��m�

ڬ�9����3����RM������0�	�ip�����_��7�D��SA����i�w�[��f-�A� r�/�'�Z5���=j��gݡ����so�mK2V��?�a=<ɱ`���ӛx�M��0��GV��g;�N\h�G��L����Qc`�T<�(�#����b�ѕ1}Cv:�����f���?��B����$�
�������}�B��Oe*-NuKHWZ�'؇H,
���o A���!�3��d����7�W_��\M*��T���O�X1�	F�p�d��-	�����i�C��̛j�1ǟ v���q���!ML5�2�����жY��d*���ȥ�^�����]8Lg����(�q&(��F�.='���.&	K�ar�0tS����x��[��,C�)}m��H�@��dr�N'�Ȇ	�?� #�"�̕�A�1k}��HVģ�x��P���%w�Z����?GGq<�(^&: =XS}&������L�H��N^k�Q��MY.sF��t�.�&����g8$�W^P�wF2!Jr�s�2��������4HM~�$�*�̀��Hr���qA�ڪ����M°Fb�dѳNң'MB����ڂzM?�'��dJ`�hk�4���U>2'"�,jr3y�g��{�3 �uA4G��0-�Ƨ� ����L��)�B��F��Ӊ��R*<Iۯ�F܍:,�b�s�̷��w�����N�������WO`�2-_]O�ݰ�C����>�T�u�z�U�٧�'B�#�#��g���z���u1���Տnmi#x�B��i��T�w��K4�D瓽�,�+;j�����د Q� i��*�Ѩ��|�A�q�.��J%��].W#Zi�y��'�;�@ߺv2=C���D����5��bO�'��P��1�BrC�n���ŕ*@T�A�y��^N6P��+u���+1A~s̪�	1���Z����jZ��"�^��f���iQx���)Z�b������[]c�D��%������\�F��I�'s�1�Mѝ��:	���i���L�u���^]�	��R�|:��}��� "3ܔ�҈�
 �^yxC��rp��� v��M\�Y�B��L0dQ��E�w�k�U���U�#��ݝ��J���-��|���q��J�!W�|�V[�_�j�5�%N�w�o�$u���Rl�Ⱦ�<�_�3�d]2�et8��ռ9��-�D��l���d��� tݱn�('$��9���~^��E��_ٚ�+���Y�,�ī��R�9Qw��L� u���9���Ә2_Je�k\$t�_�3q-.��� 3��E�!F�>{�{�Uz��[
�D�n�	�O�>�� �?	��rW4H���z�o�ߢ�͌Z�K+�8Ԓ&�ϐ���!���h�^FXB
���x_b��V��=`ybS`f�0E |�.d&	��O6�w�+�n,�s������Y{�/i|G��.Pc�Y*@כ�_%�̈v@)��W{��u ql!�� ��/U�����∲�g�NS85�y��_��+�j��U�MjfT'	Z�&�o/T�찼��k^oG�S��̊�7Z<�?w]�g/�1�4��D�|���r*�	��ʩ�a<����e�ξ<q�������- 	�a1NA�U��`�ZN��N5��<���4{Y.ݨ�I�����3�t����h�5hc��Ԥ
��e5�hx���d������`�7��Jo�+;1���ϸ��#ˏ����X�$��
�;��J��~��nN\ui���l���#)      Ĵ���	��Z�Zv�J�(��0���~"�'*<ac�ʄ��	Z,t�P���?Y�I]!5/4�95� Pv���J��S���e�Nl��?i�|rꉣ��Ja�b�ݲ2��R�`9�����O�`yڴ!�&`r��;s�Ψ�cFէ@z�Z+O~�)N&�M�BB3ΓE�^�'�T�#�)�4[��LK��ٟА�z��&�b�H�O6O�����d�r�Xp�%^�7�tM8Ue٪U�Fx�
C�'T����Uqp��x%L��§^�$��$�d�2�i�L�O�]1ҏ�<��A��#W�3�2O��؎�D���Or	���I@Jlӳ�^#fڼ!�$N�'��xDx�k�l}��]�� J�cV�<����gF&��	�D��cb��_�t��� CL�̘�PϚ2Q^�f!W^�'N,Ex2�I:#>�R�IЩ6����D�C�&p��}r�PQ�'-��'�S���H.h���.��1�*O�@@��d����'��y�f-�1d��d��kF�V�\4Ն[H�']ڌDx"�����L�>\��*'��c��� 
7�	 c����x�$ϑ'��B�#L�Xz$�R�#܈�~"I�e�'i$�Ey���Z1x����S�Pv��އ�?�M��A��W��|b������w�p�&�� j��5#%�B?(հ9��{���k�'��	�O4� U�D�Ů�ȗIđ��}	R�+��b:Q����r�:H*H�>@{B4�"OR3 �  �N���x�J6�~�B��A)��ޑ��4�c� #
<�/bKϯ�DmF���q��)7 �����9Խ�(k���z;5�%�
���^39?�-�/Ь}:\h��&�ȹ>B�|V{��_cH$����=r�	�E��,倴��*^������Y6����rÏN��k��x_/w��P)mW��J�	�(��5�*�	����+�p��EO^�q��
���d� �ߟ�5�5���iS���� ^h�-�|X�Z��o��"�p���1��b"������������hۗ&Ď���S�]�@�Ӿ�D�ad��>ډe�U�&�NRXJ�	��SS�h.*
\��2ٷ;�	���5�`\�V�n��K�@�U�qr{V�t��<.��T�8��Y1�_j���3�t �fQ��x��y�q�6���z���pʚ����ԯpUO~��d] f�9;"o6!Ɲ����,m �є8�?�D�	� �j��j�ǆP�<��D�u�'�!t�K|   A    :IZ@-�nkZ��&C�'ll\�0bLz+��AI��e���؟8E{BF�:d 2  ���������b��X[�   I   Ĵ���	��ZXKv	�+s��0���~"�ײK*<ac�ʄ��	Z�q�\x��g�R�m��NS�{���"ˬ�� h���ܴ���a����	H���Q��+�I&;t�ر�\6B;L���_G�']�Dx¬���a�S͚�ڊBv%�*r1�%D� oy��F�_�6,oڦn ��(v����Չk���:<��(qd	�(�D��G
	�$8����4�v��O�L�	��u`��?�ɯ+�J`�0S�:�ĐjsK��MƘX�Õ� �1O�������(O��a�'��T)E*B 1�vŚ�f�h �mXI>a��4�'l(�OR�yS�D3-t��cт�"���0O��Ȍ�D	6�O )�"�	6]w��c�j�$�Ԥ���~�'I�LFxb!�k}R�˒Nά���*|\<}�A�	���ɋU�DzA���;(�r"��d1ڀ�(7��j�Q�'^Dxل*�˘o(� �ˀ���}���Z�'�R��'C�9� �֍J���D��H�\+/O�4������'�(�Y�*L�R ��T�*\	R�d�'�ʬGx�˗柜�Q&ʱ&�(��SH9���Pa0��!���;T�x�	����F������Β�~��I�']�a&�,�f�FdX�� �~��ง�ÄIk���E�~re�T�����zU��c�i��xo��Q����*F�a$�g�ѳ�����&�a�	�z��郦�?񄁹�r�虑
����cb����`wh�jQ���Q�I�0��G:��!Hć�-:2�C��xN �  ��z_4�@w_��J@nN�	pXe��CǍGm�<i�搬#�t+G�L�a���+ҍe,|�I��M��i���'���'xB�'3���54���)���,�碀�8�4���Q`�	#^'0��B*��UhޑY���'D�P:S�Orc�̭;gغ���5kc21x�΋�vX�+��rc�(��$�n��O����$�H#�r�a`�&5�H�
�'�*�K�ʗb�`��N�l����
���'�0���A��x�h�CF�bb
�'Q~U���L6��`�sÅ `!T�1���+�S�TJ�>�M�b�C����3ˌ�tWўt��K���'!^tͧ^�ٛ�%�J�U	��'k
<��{ҥ��b?O&4%�[3'�`=�<�	�G"O4� +�Z��<h��$��#��/�S�'p���.�!  �#JL�B݄   A    :IZ@-�nkZ��&C�'ll\�0bLz+��AI��e���؟8E{BF�:d 2  �6Kl`
�9�<ig�   �	  �  U  �   V)   �pA���D���\�'ll\�0BLz+��A	��e�2b��UA�/Z0�'��ث Q�0�
���C�'-U�0�Gg��<PI��'_�]c2��(�x�;
^%nY6�[1)�(���'��!��́�2����=.���5d	�?�����?���'���(� �#N��pv'��6����
ߓ$��'��]���3	q�M�d��g����{�`є:�b�dޮF%��5sI�H ���ytX�����x�'1�����'b6��L~��V9VL��g�	q��طa�g�<	d�(ٌ�e��W�}Ѕ" f�� �?qh!m���[qD
x��@e�G�<AB`���p$��..�2��B��%둞�'|PD�K�6E���H�k�t=w�	(� �s�y����ʲ��ն���
�qqzUy�d����'�V$ۅ	u�g��]��f��@"���D��C�I5�<L��JP?��0��O��"alb�DE{��� ��F��3rG�|��逥혹�y�cޖ�`�j
{m��ٴn҅U����O��㟘i�N,5��
��Ϟ�E84J�O쁩$fW̓�E�ԡ� ,E��S������,[�"@ؼ�Q��&��?����!)����>�`a�-�h�<�� �$b�TQa L�4ᄨsp�b�'��y64.�q��JE�yפ$�yr.��L��$I�Ζ�DQU)��Ƕ�?��Q�X���$�g�I���rcƼF��c�I����� f�0;�r���̨[M��`��>,��v��#q��K�&��V��@����XQ��#�I#t�K��.Q�������d]xab��=se
�m��=��Ș�$@��p�/٩gԮX�u���Q����,� y*6Y�ëˤ#��$Y����R^��dŦ	�ܴ�?i��?Q��?�����iY�C�L��'^�j�J��S��'D�{�o!��L���2@�Q="e��"�qO�U����O�b��2"�.+���K�	�is#[5[O��qa&ܚ��I�}� �>�ɣ" t���j���0PJx��S	:��"Op�pb*�,J[��9�ؒʀ��'B�O�}�!O\�Z��1"k_)ZX�p�"O���u�� 51�p�k*�l(��
r���i��O9�pM��^!�g�\kU��<i�SjT�����?I*�Zq�2Er�l����Y>h2P��ܲ�>0��ߟd��$<� ���I DlҧJL<��d�$ybƤ�B��80��d�r@YF��;A#<�~�"�	T��P�ț�1}B����[�I7.����OT������J�Z�q e(2'?�ؽY���O����لq��+�­<]켊Ҏ^F�"=��O4��Rŕ6tcx�'���d�(Z.U\��	���x�'��!��֭9	�O,QGP���.K�;�X��bE�>	�JiX���T�A)f��:�)�GF�=u1�I�Dc����)<�4P�Ǭ����I͊�:q>��K>qG�۟�>O�����¡Ct}�q��4R����W"O"Ei�cR0�D��Mإ2˞Al�'T��PF�"<��/��;on�󭀯�u@�c�+I� I��$�5,��X��'��'Z2�d��I�'���ƭ+(E��o�'Y��b�-L(UU�Iر���a~2*�!���!-D�昙�G<q!(�!�E�0?�"8F��4b�#�Pf^xyv��x��ݟx��֟��'q���Ց\���h�@̫b�r���K�T��{��:���̩��/[ sڄ ��F�2�qO�m*U2O2ʓ] �����<Yٴd���%�M�R�P����Ϧs�*KV�'���Q�J��3e�'E�Ʌ$e��k%/��J��*�i>�5е�ݴE�
��#�,�˓H䜹󂁊{M��*�NJ覡â!��R�F�� -X�)L�]�R&:,O �8��'��6m�Y?��A��9\:���D�~���zA�r��?�˓(5~Y��$Z
3�x�*�/���?	��~R�ThΠB ���u����H�δ�����G�wg&m�<���$�|��*޷�M�3fѰa�(�t`�(vl}xg��5n��'�5D/B��~�H� �W��O�b8�s+ϗ��F̂���pB��
o>esǃ�|��5"�������M�B�)3�:�'��}pd��F�j���}�$��z���Ovl��H���ݘ#�0�c�лB� �"5���\ �1
�'aX�S��ݾfX:���6`� �����`�@��J�!����B`�t4���U�h(^����KR�'�r#!@��'��''"��g�? ��Z-H50�b%���P����:n� ���<ii��Od�
2�8�L<1�%�K=^y�h��h�9I� | ���a����4��p�~&�c�׽������M9ܰL�f��EU��γ<ٶ���S�?��>Q��F�f�6�15��z���i6�E�<Q�<碐�򬍛m�Z}�C�b2 ���D�*gx�@�����D�s�tqu�ןU�(AZ���o��$D�+A Q���DċQ� �Pa�|B�-pc�%����r����J2�y��5�t��A�}���"I��y��/�l���|z�)2�[:r���$+I��� �"��Q-�c��{&!���HG���2�Ϡ� �pb ���OZ�Gz��/e?����	�u�֫��b��I�aI�.3��[>��ԫAH�B�e&?)i�`_)e���:0K�&����8D��q�IP#� ���T�� l8LOl�(h'������
oE��(X*� 6D� :��6W�� :��"T���K)8�ɣ�HO�S�,y.aR�$΁=/B}b�(�kҘ�*��F+Ch���<����?���pBJ��C���Tp��q̓:*�ur&?�3����y��\P�@�v��PMԧ,�!�D�KRU�At9�m{A[K1O��=�|
gJ
��}k�$�
"Yi��M�Q�<� gͣ=!��a޾Vb���j��HOR�'��Of8�.�;v:���E��3�ҭ1�'k�	�Tb�(����`o��1�C:u�E	6���h�R�/Щ&q:�����\��3�
�W�V���B�e�!�d�:sT����i�8V�h�@��_��`��ɤB��PC��Ö)6���#Yg��C�"�~�
g+L_�����a���$�N}��9ғ4��'̀�k$<+�PX��̰b���1�'q�T�o��'��|Y����~D�P��<�\�2��.d��<�ȓ-e��%/�8AA����K�6�����:���1I[1"Ƭ�"P7���'F:�q�O�.0��2�E�<�l	ߓr��'�$	��T"p�YB�~,���G?�x��I��'8dp�� ��|�Ef^%�(�K��9�*�<X�0c��cQ�=��-dN�I녠�4�]t*ݸ�*JQ�<����:H2i�Ϗ,8��}H���E��d�?�ģإ:��1	a�E#u�d�A��W�<�%C�(9H�0K��"E��u0dhT�F���'mb�����H����h� K�9��I�7y��	�y�0�"6k(L ����Z�m�����'�h3���d�g�I�>]Q�'A;�ȋcK��	�C䉘Bȡ�EcI���H��.i��:�Ş#�Z���P��F�k�<{�J�<��5|��B�
"d	4�	�O��HO�ʧ?!�OJ�ʒ�H$`�FH:VJ�#Z� e�'ێ���;��l܎"|ڱ� Sn��n�&5�|iK4� J���G.����>tw��&V�Q�!�d����]X�ʞ�N�P�Q֥W\]����I�`m�E i,9��ЂfeV,tC䉖hS�)��J�6�XZ چ*�ĊM}b(=��'�\�s����:�	s����'&xl�!�ۘ''��� ��E�>����E0iN}SS�N2y�!�ȓUԅB���#%@����N-P�:m��0dT��
�
n�t��l�va�
�'u��(	�4��h*U+߰dز�!�5�'~J��V�	�P�f!��%/_����	(P�t�	��N���'�.v�����x5���O��%���1O����t,��cT�3&"�I�)K��y�jU�,<D9)`���F.��x�R��0=1�2���,��e��@ ;��� ���y��6q�<��	�+�
��w@���'��"=�O��ɑSJ^8+h�� �.�
$�ґـG"ғ~�5���|��d�38CJq��� KԽ:��T�h�1O�@3f��9����S�? $�x��wn������
��M�U"O�)�k��U;R�yх[�&�\m���+�Şy�U[�� �h����M��	!�q��{�J��C���-�v��4��#�򵹋��|�C��pŉD �2\��@��W�r�#7�^b�|0t�Ӈ<��Q���]�Gø�K��ms����[
�����ɧ1Nh�iB��%e���&Հ}s�C�Io8^�9bF[{�����2e�v#<A
ϓc!����Ev X�g��!e^�!�ȓGH��YV�0up�!�ʛwq���;��D�f�'B1O�����kg���vjG�`>�L*��O��Df�,�1O\)SflE�'�Dt����:���"b�]��i��'�ּ���څ��iҨݰ!��z�'4N�P��U� �j Q엍4Z���OR�;��/<���Ѱ@�>�z�'��OP����j��BNϙv�LX�1�$0� &�	cu�'5\L𶭉~�(��$3�<��J���q�4�Hb�8�U�3�	Z�ט%8�bG��4#��KM"!��6-b�`��r� M�Vzaz"���W��j'��q͌�P��װK�!�Ğ�K�f��܋�@�x���6^o�O�Dzʟ�E��+�Mt;CȌ�a+qA��K�'#�	�`0�I+Z"�.�$f�P}��*����cǨ��Qdb��q〝��q��'j���̎��ʱy͏&y�x�)�'�\ r`H�!Ј0ȶ	�o���y��)�#Ni�˃*�x$�{utC��zo�J�F�'0rm��i�YtPFz�Z>����6���R�R�R�8�c�B���?i'��11O��`��c�~LX��F}������9s�49g��|n���\9O�4�	=Up��$�N�70!�d�����g--f����an�@����ɩX���s��$L�&��q�F'zfRC�	�=Q�Jvꃃ+Z�Ȥ@�����A}��*ғ9��'���pdH�AG��%Λ��ġ�'�H�9�`���'�J�1�@���]5�5a�� /�,�e�O�R���'"����O�#٘���F�K�8P�ȓY	6�C%¢8Ό�zp��/`�^��	�'"<��mV�>/� (�\\J�
ߓ��'Ǿ��5�98 E��L�'�Xb���
p�����%�dݲd�T� ��&Ō���$��K�M��_�1O@�I��d���ukZY\<��v(-�y��@w��M[1�=}��-��A݇�0=a�B�O�f�|�$�ĩJ�V���,�y���7\(<Y��CN�q���'��#=�O|v��AN��&�88�F� � 1�8ғY8$$�P�����D��f�D �vb�A��eگyLc�D�M�/9�q��'� PƨE�I��)H���3p6~���'�`�	Kz����[&X�ْ�y��)�S�M�j}Z�	�>Ũ`С�ׇ#��B�ɤ@��r���2#-�(��MV%�EDz�P>uY�"�ԚJ,Jю�3J&���!�?��Nk1OL�S�6
T�$��DU�����ХB�l���6B�1T��DN�"�t��|N�I�ŏ���!�䋚76��L��T1N]��.ۦ`��d��I	B�P"P�K7X�~�Tg\�]|>C�	�h�qT��3XL!�$���e 2��HG}b"9�S��'�Zͳ��6X|�����ax��'hN��)���'����)��y�d*b��?r�kGC	�$���ȓ}��xv����ܕi@�E$jD��`k���d�h���9�b�QT��
�'�,��-_�Ze+��Y�uw^�Cߓrm�'�bܻt�_��|:¬(E��A��`<ғEFM�0�'���+��}�q�,Z���QReDK�2Vb�0�� 5���~۞E�*B�3:Abr��N�!�� $�+@�]�(�����䉠xd����'��O�\�(I6-i,�($��4���3"OZT���Nu�1����cԞT ���s���铿7��p��9.~�t/�3sd�=���<91O@͓�O����1��%A�R9A��+v]0l�0��6�0l���L>96�_4E�ִ��kM�QĂ�_�<���
	C@�-�FƐ�M?�l�$b�b̓�hO1�\H��(�$#�vUs�F
_.�(��"O���)&x쳵�U�p<0=q�.ғ���o�4
�T�ӈE.l�h(2��pd��I�9r�9�y��_e��?1�l�Ma��""Y�v��B�\s�V���1�*�j�,:���r���P
Tl�ȓa�6����F��y����5Td�Fx��'�9�.��v� \S�Cl�z���'��1A6_�,�$`Αg�`��Z��I�HO"c���懈�2ܘ �&��U��Iqv �����4!��$Gyb�_R�,Ol*S�qBAnI�RJ� ��i>D��!��\�(�FI�E�2�q�?D�Dc2à'y��3ЫQ$` ��B�YTh<�g�X 9l,t��+�$_�0�Fl��lCN>1�oF�>��&.�7���!G�Q���hO�n�\���W�$�����o}:P"V����'��<�&�K�ӆ�L YqiG��L�+��L��C�ɋ^]n`kD
U�����ȃE����;�I��\�`�S�E���9�O�12�C��(v�hM+A#_��%����`����ь��?�h�h\�0]�9C"fӏY�ΌcFl�k�'.�����3�	�e.�)Έ#��� ��c^T;,���c�T9$�TEq��'�v��5�C�v��T0��I� �q�'릉����/ d�MJuΊ$�`��yr�)擵!B<��>�D�bb$SZC��/A5���-� ��kc���Dz�P>Ţ�� @�@�$��(y�Z@����?	��^�1O%���'�,���%�4T0 �C��KZ�xS�Â����G�d� 唳Fϰ�+$�I��y�1p*�2gnޏ;��々��O��$Y�~k,u;�,߀1:�Kr�H<'A!�mdb5+�$ ,¬�  �I?B.�>a�	K�|A�0��)t	H�"�O&2s�d��q~�fO^�(O�cI>���Њ��P��x�T��b�<���Q7�m$h��ѣb�U�<qį�EЎ�����خD� ����xR�K(�2<1�0Z�Di��Ȓ��=�!�|�Fќyl��<CE�I�r�]&��'�ў֝3�*�$E1&qIR����`!c�\�V�Oș0�y")Q'��'@?�JÊD(�(�0V�V�[����ȓ*D68��JȰu�H-��M&P�\����Z��jݘ%	Q�T���z4���(��}{�A�� F7k0��Qԍ��kJP�?�s�)��.A�wD�#��8 y��2'딋�hO�g�n̓���?I����$X
*E��X0�U�R����<Y4�E�R��>�O�%��b�5�e+� ��z�2�T"O
�ZZ�=҅H�k������_ߘ'yўb>ţ�A-&��Eٔ)F
F��)e�7D�$��oE�.^(P��C�ξ�x�BB�'��%��'�����L{:0{@l��nQ�]E0C��A�(�"͆	kl���}��k�"�)Rl����'��� �g����Wo�6(�D���'*�hvF�R�.�Prb�m�J1���-<OX|��O��F�Hs�!�j�5D��X�α��5	��*{�a@u��O��'pV"=��yR�C<0����O ��)tA=�~�����剿+��'�"<����?P���6f�3G �A��'��d
��3��5��O-<������ ��8���.\�tD��o���V-��84�PK�;P�v�	?�����/|O��&��A��&�p0���%y
�5��#�	]��u��9�?Y$��DdQ%�
�6��L��̘M�v�nb�ȫ�=�ɘ	�r��jNzǔu�D�5;�!��b�l96��F�ȹp5+D��azB���>s�`��'�N�˅P�!�Ĉ��1��\
lY,D	�O�,EzʟR8	g��4/r��C�L�_%F�"�2�
N<���$� ��D�"nz��q	�0/�X��H�
vd1OX��@�*����&�ذ℄%B#2�P���݆ȓ�`���R�N�9���]�C�j��<������`���dO^>U� �,�=,!��(f�NX�A,�;)��y���Sf�"=1/��D�?IM �/Bѻ���v�R��Vk��:P�����d�'S�=KEp��I�OH�d�O7���_L�9���
4�1�ת�i"��A����l�
�����ēF��iG�Ð>��dҶ�	�!Gđj5�-P%��'��p�H9�3�щR���0���+����7e�f�U�IC~B
��?ͧ�HOBY�����t�`E�7�U�}8J��C"ODuц�Ãa�2�S�B��P:P)*=O��I�:+�"<�Ӝ�?��O����ˇ!J�I�$��*���tI;T��6�6�O�yk��q��lA�������Eɟ,���&
Þ�d]�퉈�ڥ�ɑ�H����GǞ�V�ɔ��1���%)���=	6�+I�=h�L;Wjf�5h�^0 -�IϟdG{����a��řOX�q����D��\!�$5ChP����'���ф)�X�qO��d��O�˓7�� D���T�i	��9�E}<��#�7;B�����Oz��?y����Ԣ@��h���
M
إ�2!��$�ٚr���*,(D��a�����ɍufx��F�%΄�+1JH�B��I(��d �<!��-"t�X��'7��I��'3��@�S�V�@�k@c��*� (�{B�'����W�A����$`��$������.�Sℌ_�@�`8�u�� D� �ĥŴ�� ���V�r�td��?��d;�_w���gZ�m�&� ��ȷU$�Y������d�O�0BV�ϝ#����p�-_�:i�i>mXq�B�~�� �T����,z�&���>��p�d�1R'�O��0G�(�X�YMܜ5(��R��?h,P���x� ��?���h��69&�Z,V�m~
��`(�i����ē���1I�W�
U%A��嶵��	��(O��BMȺ��)���t��zpkȉ�MS��?A��q���Ӧ����x��|}rEB�#�ּa�̙8� 2Wd�/_w�;��q�N
ڴm�n��&��D�g�=W�� h��'�D�A4'C�y,^YV�Xb�
�1�mk�@�y�	�p�g��4Z����0/�%@qpx@�$pdM�������"I�OR��Z'��4�I	('D��gI��!�$M�������i܉y��,j��B,����؟��'�L)�K]�Gt}#`c�����$�L*	�ְn��L�	͟ܕ'�2�'T�)_��n�K�ܘh ~���H�w��ͩB
���$Je؞ �7GT���[׭�<�X��#�L�?�Y�CB�e�(t�
ۓV9��Cƙ,�b��Ń�yx4=��PʟT��U�'Q�O� H�@��?vSRK2W@�"O�Ȱ1f4t�0�aH��k���PU�$ʦ���J�gU�l�+g�U�pȏ��`�D 2p��C䉎G�˵��?k�Ґ(Ŋ >1VC��l��E�î^�ʈS"Iݎ
��C�	"8�"|c!�#�t��q��7��C��9,dB�h�-U��e�E(�/-l\B�	Q�2H�� ��d��5`��h0�>���\{�O�ldb�� ��M����9	�'���I�9ci2L�qNЇ'2���'&JK���t�j�	�~�ڥ��' ^�h�SPÒ��Q�F�s^��'��LG�Θ7�9@�^�=�X��'>2�#5 e�Ĥ�G��=�T̊�'H��� ��    i  K    Z  �#  �)  /+   Ĵ���	����Z�,C�'ll\�0�|r�'~i*���i��� B^(v��8�'���q��+�E��oE��.����qf�a1�r�~X�m��!阽q�D9����m@��~zS�m����q��l;�\0�A�(Qz]@n�$S�A�u�Y�ݲ�$Բ�N@(��@c<qC�"y*���m�8r�ȓ�_�g�v�*�-ݐ� D�#�A� @�Y�G� �Ov 8Wǔ�u'���D#�m�	�"O>	W	NS�q���B�Q8#!�$e¬���A?���+
�>!�#S��ep��_,K��2p��!iG!�$���t�BA`�qh��i%)T3B!�JH1t9�C숊]e�M����'�!�d�`16ik��/Xrڵ����!Dg!�$J7,��r� V
W��X0���$Y!�� V&]Y�Ύ����
�ex!�dC϶i��G�M�������!�ć�C����@��q���ƍڿI�!�$��S"@��UHK|j��ѫ�!�$�<t<�aI�K�[CR��Ӄ�<�!�[�z� ,��X�!�0���'W!�DD�'�)HE�L7)�Ny�5�Q�4�!��u��騣�\�l�t\���-/�!�DN�Ix��K� ����ےV�!���R�hA��6s�b�[�dߣX!�DC!:�(��N�b����ԥ�g�!��2�����Ҫ�br��5�!�䉱[�
u+Ʃ�/皅c�/��Q�!�$RM��0��=l��������!���<!Zě�B��ay�!6R[!�Ě�n�H��%��u<�U���Y�!�d�6�"�I�%�/$�j��5�!�������	X��}�Ԇ,P�!�D�7"p�B �P��AA ��/0�!�D�8�`�§��	]�d�'k�W�!�$)}(9��e�3'�.��U�]B�!�џ�V�a2�@)i�X4�AA�z:!�;ƌ��D��Uܤ�E�O4Ha~�#4",��0�@Q`�`�2ȟ�n�I�M,N�E 4�		3 �8��>lO�q�+�w+�E��K�.�b��	� ����jͪH^�`h�U�al�7�����䎒{[�y!A윊��
G�<yeoY-��4K�x�bU�����<1�f�?k�Dف�.^5y�xhzgkQ֦#}*!��-�N������\�������N�<90.�0�fa�ɇ� ���7���c����o���� K�6��1�̟�t�>�'�/<o���Ʈ�5��|��&��tj��.I��Hx�O�<��x�¨���������w9��p󬅷�
@j
��ιyb���p@�/�>�nE|���)}��	ch|� ���M��Fg�U�.��J�������Նȓi@><�p�lS*�2�LW+F�U̓,���4��;C��d�U�I �<o:ҧ�89��(
R�zED��Z�Єȓ[�E�'!E�n��i�ʛ9f>���HX\R�lZ#M��y2��_�����v�W�1ԌթG��M�H �#1"��Ɂ8������@�ܔ�T`:���&_�3Vf�
��U)kEf���Pذ=pl=�]�B��75h�-r���E�'C� ��ߏ��
��%����6�p�J�Μ�NH���jޅ�+#|jB�&��$�%�Ǚk�d`�O�F�I�|������Y�`6́��f�nD%ɏ��I%1Mh�8���N��p
�`�(�!�d
�z~<��N7�	��4&qY��ߓY��p��0�8B՝?�(�}�`B�5i�4q!�K�sm ����\��0?�C��g�ҭ:R6_cv�Z�N�9	0N۟c���b��G(���'v��X�(�?D�H�
G��Zp^�c���Ʀ~�$����;!��1E�;lm�;N��I�0(�(y�Ek�"�.����ȓ8̘	��"�y��\�5�)Z~�Eϓ
�y��#յ;�X���D�X�����X�Qv��<� AKG;�@B��8+�\�8P�ӭ�B1VK\�N9���T��c���H%� uD��!���$Z?`�tp�X���� .wa~�xيЃh�? �ARc�@�gU�D�hh�h�,D�v�HY�Д��I�N��ᕇWy���# �U�k�#>����R|r�'��Ġ�	ra��l��N\��\��b�:z�a��>��L�ȓc(R��S�����a�?$�~i̓n������S����@�㏶�ҵo:ҧD�>5�����#�!��D��|��,晣C� �J��I ���"}����n�	Z��nZ,iDt��G�׎���s�~P��T������:%8l����2\��n���!Ԍ�6R@:��a��	�aR�c�-"h ����=)�/ͪ= �@ⰇJ:C�H���Mw�'%x�X��#(�vQJa$91�:�����k��Jw"�24��/0�x��D�q�<�0/� ��0�)Ŷ��!��_L�ɖT�#��Ol>IY6fG ���b�~�@0�@#D�t���J���0�K��9��P0��R��'ƸXD�,O����F#*���#<IUV�0�"O$J0O��.�|)���y(���"O�-��L�,05D���F�B)f �"O����Ⱥ��|i�ꜳ]{p�*�"O0�aqFX#Ty8�P�B;pPh�"O��I�T2��ItN��{���H�"O�xCD��0�DYP��Q���1�"O@�V@��(vJ��@�͖'I��H�"ON����jv�YN�c����"Of��Qo��v:.HKÍNH��P�"Ohe�կՔ$����ǒ7@�V�`"O���6�\��%�ƦcC`�J�"O %ÖƗ4���哆~�>!�"Oj�8���1t��ukNS�Ȥ��"Oj�ˑQ�rD����@�TY#"O�iB�"� '���kG������5"O����	�#n�v�Y��Xe�aۄ"OR%�ciJ�fM�2ǣV�}b88�"OĽ1��*<��A� ��{.�$x"O�,�cA�4J�(�g��7�yZ�"OjI9%BЈF�\��"��1��"O����ɮ3���f�.� �1"O����� q	��	����)��KR"OXd ���^v&�PF�+�,͸�"O�� 'c�E�:Y�@*̤_d*q�"Ohm�K�E66p!���,B�4�h�"O6�9��zZ��!�1	.\���"O�5��2Y��pa��3��,�c"O%@���<ZG�Z堁�Q"ÒHd��-~hQšҮ̶�1��'v�b�]��8'H�/�Fa�/�#t�X<a��3D��0g���t2��w�HP)r�3�	RԊ�o�|�O�V �.B�h�"��j�{���'�t� A�<D���H�o������ B)R��A S���/2�g~�i�8L�2C	G�UCV����y��Q���c��Z .M�c@��z~D��B�&�@h��'T�Iad��V�ʝp�AĘ\��C�->�9���q9�8���i��%pA'~�2e Fd*M�jx��"O�qqX=��hZU�<M�f�r�x��78�� �� r�� 	���_��"���x`�`�4T��H{�"On�{U�� L��C��+!�Z����� ^Sz���B����t�}&�hj�LF�����*
�7ڢ���-�4{"k�6_.=#���s��{2M�� W�l����b�(�8#A�gSaz"e�%bŸ�ɔΞ�T5P� ߆�0<)­\�4v��
���2Gx6�6� " ��͓ G���&A
%2-���'J
��;9=ҙrW������W~~�+�	7��H���<�J��y��L�!�[3V�J5XG�M0T����"Oz� �
�2s#�l*�¹;c�j���.@(�,13�ۆ�(��7�݀V�1�(�O���0��y|�`*�H J����O���4g�B��	S@� �b&�V".D�0*���E4Q)b
�)������&@iB��� �̰��OF�ax̴5$"a���U��1�ac�� ��3k�R�*@���C�b�cJ?4��x��WH��X�N���3��,}�f�t�~bcL�9U�0���U�Ovĵ#EM�V�$;၇#���@�'#Hu C��>s��!��DQ�j0�D'rJ�1c�
"[J��M��Ƹ��
B@͉��Qa��0� ��+�P<�ȓ+� �6`�m����I�n� ��	0/�&��bB	=9���D3g>���Ѳ*K��Q��3.ka{Rm��j�`�m�0d������l8M��cR>�P��vD-D�pX ���J��a#�-�T�1�,�I+zUl1�i�>��>I���m���AA܏KZ~8�C'D��w�ȯi���F�
@H��B�07������y~��D����V� qA.`��`��,,b!�$�8mǴ�y���7C�`�� �^Y��制yotP��'�@t� �_ �P4(�$�#6i�� �e��K/O���뉋N�H�	�g�ʒ"O��:���.=:�Y!���#Ah�"O`S��؈U�L�ɴ&՝Þ�B4"O���f�އ�f����X1�<�"O-�"���5Y��%%��?u��"O�ͫ��i)�[g.V2Tk<E�#"O��I��0��c�� �*ȹB�K�!�d�"��pD����4��l׮{!�*v�3a/��҈Ӈ�5p�!�DF�0>-�B� ��݃ECH��!��42>��b+�#s�����AżO.!�uN2xB�m�1�0m�j�0!�۸���E�U�L��CO!�PO��qe�_�D2�����ay!��} ճG"g�$TĚ:�NՅ�v������� ��=��?Zԅ�����C�Z�R��U�5m�<��ȓw ���p�"9B֙��	1|�r���o�V��d�M+%�\C @�	V�����M�1�$DF9l
�����L�ip�]��uӈ��f��K'�� %X�/�<-�ȓRf@�Z��!	`%�pÇ))�l��`ՠ,�bN^�(*,*s�֕ԑ��C� �c
Q�1r�K�b�*����Cht�`E�	�u�C7c�-�ȓmoJUH��ʸ��̇�R��)��u$�( k�J�� �kJ�W=^]��O� �صe��()6i�Bb��^<�ȓ%���9W�&��dH� �
���ȓ�TP�U#I�d�H�x��`l��ȓ9\v��Taƾ9b�h�K��5�����j<J�@��8�h�NIv(�ȓ3��tꦬׇ&����2Ót��B�I�����"H�:&��)�V0��B�	�QU�9:r!��6�LY0��:PC�I.N�4�����'H���dF�h�`B�����p#�t=���s�O9n��C�	�r�d��ԍ�w�� G�L�^e�C�$n�Żv+òU\(��@�5)EC�	]UF��v⛂DU�h� [E�C䉨 &Z�@�f�*J_����>X�C�	��8 �bI�>�*(1��9�(B�I�;�DM�S&FM��(�A� W
�C䉑sڈ	a,��#�4$p2fQ+e�tB�ae��hg��L��1eg�$DC��8c]�����\�c�����C�[ C�	.Ty�Y��i��(K��%�)t��B�4]�Ă�ć>|^`b4�B4}=lC�&5o�K�(8K�x�󁕎)�<C�	<���.
�TdN��qnw�,C�)� ���jF+J>���1�	�+u��"O<LR3��;��rs��N�h�"O"�)��CĂh4x�q�"O�I��gZ����	sC����xR"O��0#�;
�t���}un��"O���BM��i�X9��12C\D�d"Ohs��;{�$Q�"�'�Bف"Ovu�Q!݃Z�LQzT!' �d-��"O�䐗OӖ"���*��B�����DY��m(`�TX�`�G��^��i�&|I��� D���`�ʖG����[=t����$D�#���,�cdE�"7 �EG6D�8ˆ�����X���<%L�[w�8D���I�4�|Lz4AS8 ҽ��7D��s2�$"���'B�D��9���(D��Z�]�~"n`�G�U �˄�&D���V��@A�|"�
�3}���(2D�|��쒰h�,#w冴t�H� ��"D��(�f�r-"X�aFĽV�D�3Q."D�����>0�RE���I�
X��%D�$rr�מ#**ua��ުv�tY�8D�x�FA �2Lx�AC�fh�15D����^dht8�V�P�B����d�4D��u)�
�΄���)�xP �1D�5{�i0C�^�k���Y�!=D��e�ǒAj��[� �P<D��#Ā�O�y��K^�~vIg�5D��r��*����[�U��Еc6D�0xFG�\���g[�k%J!0�*/D�<2g�D� V	�tt4b�!^�<�c
;!�by�G�T�HB��ZN�<��F@�}(���鉓x5pzĉ�I�<�*xRh1�B����g�@D�<���.'(.�;I��{r�a��I�<i�� W�N�y��!w�$���g�x�<a�G�K���F� � :ǩt�<��-��)Y�cUkH	y��%�m�<!0��J�T8�B�,����Ac�<Q�&�X�`�$0�v����`�<)��R�& *S�Az�X����D�<�3Z@|��fƗ?]����k�<��زE�Ti#��(�N�\�<Y���!	�2��C�B�!��W�<�s�H='L �0!�
D5�Yq�MJ�<����h�Q�)7��E�,�E�<��,A�֙`U��?H�p� B�x�<��h_&�2�(��7\$l�Ǚh�<Q��љQ:b��W�+Q��
�@5T��+$�N,��A�V��_:���	2D��xs	ck|U�&D�B��E��A+D�����O��i�OC0,�	�Eb'D����Y-]�I`���+�.�K��$D��{�nݼG�đ�%LA.�*i0c D���%?����s�޺5�"!#A�0D�Tǁ	8((>P1�`A&S� %;�L.D�<�˙�J��XZ%�[�9y&e���-D�Tc�HW!�ND(` n���	h9D��� J;U�����S%@x��3@�:D�,@c�,��"h�}���q�7D��!lJ�]$.���C̹lH��kC�7D� K��Ǔ� ����F(r4��!�$4D�$Hh��J	S�iC�Y��e��0D���P)QČ�JBl.9���`��:D�0�e�/�$i7C�r�峦f-D�� H�H'�U�4.�pXW�1�x �"OL]C�+ �r'�\�0�pc"O�5�%H��" ���%|�[`"O&��&��ItDQ�p%���1,V�<y0d�N?��IV$�Z��+�L�<���+2 >����ߕe���X���\�<�gYB�<u�ë�@Y�TB
@�<��f߫A(�$l�G߮����r�<)�H�+1u<��6�\=���o�<��`03���Ɖ>��p���[C�<�1�\]��"gn��g�|�ku��I�<�E�	��0d���*{W�(�G�VI�<�U'7�8@/R�X�Ĥp��C�<�Sa��B��a���F=��U�6�P~�<Q��<&?�uX�Q�`X�L@{�<9�|�hCG��~$�&�o�<	TkF�l�Ƅ��]!XHKT��Q�<���λ�v���)>b8(�qDC�<!G��~6]�0�'c�(�IPG�X�<���$q���Z7a�"'.����(�i�<��Ȃ,
��!���3y�Rh�ab�<�bM��R6d�A����8N<QJ��X\�<Y�N͞v��8���͖;d�5NLU�<q�@�4�Z�Ҁ��)�,�"JZO�<��.��_9vYc�R<!�����BK�<q����D�1pb���&��<��]A�<�WH	�J��z�̈́3����{�<�����m�Z�{���}�����Tv�<���j.Lu��(�F��w�p�<��(�FgX�YE�B��Ԉ\E!�V�l��bs���?լ�*�݊[!��G��@���U�b5K>X+!�_ub�髂Ȟ�ύc��.?LB�	�rXD�c�)�:|�JA�͌��B�	�mL���Ǭ�5�80
�Q.�C�ɿ�v���@V�!�Y��fb	��'ńd�-�?8��Ѐ
ЬU��Q��'0P�D1)nl�GH�$�$)	�'f4y�7j<mʬ��a�7m� (�'����Ï�3Q��Y;�Tf�)0
�'�Y�$�4�¹���$[�J��	����O���Rc�֝k�.-@�ӳ�y�j�+u,���Q�A�`4�Y�w�X5�y���I8�3�m�lHP���կ�yB�����2v�N;gC�ŋ'�P��yF~���JA�fUb͡�T��y"��2�p!ʂHح�JX�eHW�yBH�]����e\)��mJ��֚�y��J�E��6.A�xl�뗦J��y�$vr}Бa�&ꨥ����y"$��skZ\��'�l$�ѢF���yB`޹#K�8[@��m����&I(�y"푀��8 ���%:�H� �y�抒�`��N�70+�=��i�%�y�+P:�p5�Wf�"
��5b��y�[+w���s��ņR^��I�*Z��y�Q�u�`đ�<�a�f�yb�I�;p�D�I\?����B�+�y�D������C�UڠҀ��y"�-Kn�t��Y�6�G�&�y��Z�Vx@��J�U}Nys'�^�y��5*X���g��S�%�fA���y+y�d�,!{����DeV��yB)��C�
GzD�`!�+[:�y
� 2(��N5��lb��@4>���"O��Y�|�D��1�@�G� ��"O ����3�V�
6(�x	�*�"O��H����o���u��Wb�{�"O� �o�J�*�4Ox�X�f"O���B��F�.0�6o�*E�ڬ��"O�h�^�"/$0�A�V=_ <;%"O��I���
��,�-�V�B�X"Oh��	�	b8]��l��Z��h2"O�	�1*F)R@0�؄����ĉa1"O��Qg�K+][�ӡ���lX� "OT�1���V� �@��L�T��Z�"O ͚�	�bgE_Lyr� 6"OT8H��S WL���T� >|s:��S"OT� q�[�=�L @uj_bj�X��"O葊胳7�H�(0_�)��"O:�K��8��UPG�#PNȈH�"O����X�i��m��GX�a$"O�9�B%��2�D�B�d��g���'"O}�`l�b!xxX�,�+h/�<'"O�X[d�Z��QI�H.c'h�"O��钧O�M�Й��́�a"f�"O^U�U�ض:.F��!J)�\��"O�驣���yհ��6oR<Vj��"Ov�i�
q�p$1����/��$�D"O�]ӥ�~��E*�m�9~�����"O6����3EE`� ѩ1qVY�"ON, �+{�PPi��^\�8I�"Oxň�	�Tof����Ą;�D%�!"O��`��`�$X����0[�"O�A�R�q.|�b��DΠ]2�"O.Tp�ȟ�[X��enJ�y��q�A"O��Se����3m �~gT���"On�ѕG�o�0�7JA1��$C�"O����;�`(�Ҋc}���R"OJ В`��nZt��  mD*��B"O�Q'�̿'�,� ]��4s�C�yr�;?��B�E9r��3�b٨�y��X�#���we�5d+`T"q�N.�y2�N�8ۡIWlt�2 ��'�y��Q�6�R�1p!K�x�1�V��)�y�c�v��I0��wb���5�C��y��C�M-�����.k�� ����y�j\8r��G�@�e��x8s�2�yB-��ԩxf�_� p#6`��y�/�>E4��AB���P������ymM,T81%kN�D�`�HEI���y�E�Pv�0���bD�{�Ή�y�9n~�{2��p�4����y�)
�}@�mʠ�l(W�]��y"P*Z��h9��K o�e�í
��yB�%b$��N�c(v�iㄓ��y"OS=S��3�#Z׾-JS_��yR,�5�*�d�T�R�~H!��H��y2 �K�
��ҚI{"�s�΢�y�)�#N�Zcn�A�Fd��X�y��� ��5����8����9�y��ͤk��*Fo�)ݢ�:u���y���3��k7�H�%В�ԩ	�y�̅�W1���V�,L���J���y�c�<$��!�q�\,�@�S��y�� 2.� ���W 7t�y�S�y��>2����f��*�Ȩ᱇^�yR��/$t�P�!�)���jR�y
� �e�Gֺ'�$s��Q
t�dl��"O�R��շ+1|�ے
G��F��"Ob�rL\	7|�樀�Me)��"O�ݚA�)��aF"ΤLmR=B0"O��
O�7�t�p�A�HQ��#$"O��y�������q T'Z
�ڦ"O��K�<;�1"�%G.i��'�2E�U�Υ?�,%���ݼ)~��'��x�0eȋh���C�'�"��'��]���c}�l���G2ݙ�'�lT���%�R�)$NI�Ch(I�'�d�pF
�o���ˣ逯Ak&��
�'�H���$� �`���Q��
�'��Y @ ����`B�e�=��ǀF�I/(ڪT�ԯ�>HE (@g�M� �C�	/�@���w��aFD�C�I�Y���k �2`�0�1��Bi�C�	�&�B�C<F��m	���LF|C�I,<~,i�(�.x�\;C�ˌB�NC�	��jM��#�.���;�HC�	�1gjY�d �N����a��LC�	~��E#�-�19��xbt�B�A�tC�	� ��5*燫`����!M�C��<��A�'j� ђ��DF�W�:C�	C��8��N9Ԑ���Ƀ�2C�M��c���8$�}2C�	�C�	KҀ���Ij��*+�?��B�)� �QiC�B�XlʲeN6:�"�S�"O !���|j��(�jʉ{BҤ�c"OhШ�E�Le*��m3z�"O�P2td��Z� �"G�_1Lj"O�aa6l
�;@�
rB0�q"OF��L��Δx�0�W�m�b銆"O��6�oD�Ұ��[��}�t"O�PPnH����Ζ�'���@"O�@��Q	[|���`�yc"O DL�Ql��pޑ�[�"O2ٸt�Ƒs���JѯC�-�`�"Oʽ���G�%�e���$+2�Ԛ�"Oz�'��I���GkR@�Q"O��2��'i�x�&�E%L)"O��q�kW7J��Q��b��`P}�"O�P��$��z�
�)����
&TDKq"O
�����9Ș���	k-h��"O���kٌm��#��e9""O� ��nB'5A��o�/5���"O8���ǟ�!��$� ���L���00"Oq�1�ƙ���}�E��"O��z5��9���t�_�C�����"O�9�Qe �p��eK"l�0Y��V"O����'�+?x�y�� �1�&�J�"O64�1�ͮK�l���b�Ƚۑ"O�DRr�S��$G3l��I�(�)�!�/�V��(�0���	hÿ}y!�ę�G��j)����f�ٍx!�E�T��+a
̝K��E��W�!�$ܦ�"-�`
�h��ᓕe�K�!�L;��$a��O�jL�9�%̱�!��Q�b�p���V0x�"gDI�!��Y�9	�90A3⏅V�!���9"-!���0<�K"� H�!��9*�ɣ�\5"�� ����!�$ݣmJ�	��˙w��d���G�jd!���if<ѐ%�� g���2*N�>Z!�$�\M��E@��n�V��5��1dG!��e�V�ȃ�I.$�
h�al@V;!�D������"W�ER��K S!�D�w�����C*awԭ�1��!���%+�%�@�vn�@Q(�&�!���JO8���F�\��f�2�!�ɸO��c�A ��R��kΆd�!�/Aj��ࢃ/[�h�a@؅?�!�G�E�8��ȑ&N���6�T�5�!��K8_@lxx�&�x����,�)�!������K�j�,9F,-$}!�� z��d��']N PH���F>!�ܦ_l�%��HN�M����K:�!�DH2x�JE�/x~4�)��J�!��>K�d囀�G�m8�����!�DȰB��e(C�L�R��5�B�
�!����P��T�MD�k�e��n!��K�b�`MZw��%-�@�E�{T!��S.6��PhA�,�Υ
s�W2\K!�$A����1���M�f�YB�D!!�DE94]�1��(̲�^��BF_!��ʿld��b�P(�6�7@J�y�!��D~Ma'��~	���o�4}�!�d̖C�.���,M�"�􌨃N")�!�D�q��D�����Ly����Θp�!�D��t�P���뀪k̄Q�ɔ 3!�F�+��X���cN!�&C�0|!�� z�h ��h)���>0Gd��c"O����f�@jBP���r�P�"O�Rf��AAX�*�d/P��l��"OZM2�k֔.��Dk0�G��
u"O,4�PJ��&l�x�c����Lac"O��,9K��M3�["4ܚx�"O�ћ���iE� A�K/i�>��&"O����IшL�TM�#���ʖ0�r"O�t�d���oVh#���K�z��"O40��+��&ШIј�:�"O8��*ȄX켸 �'猰ZE"OR�� `C��r�@ܲ_夽IC"O�5Y�����|��ċj͂ r�"O٘Ec�&���g�W��KC"O�m���m���á��3'��q�"O��a%jN�G�B�鑧�6��#�"O*�Y%�"|QЀ���N�����"O�(�B�XZ<J��ƒ0�pq�"O�ё�R^���w��/D���""OT"��:;�ra!��8dc5"Ob5�ЈɩB� ��S(KH��"O<a(�� AFPyp$��6���a"O8����p�Z�q�z���c&"ONЫ��+G��%���z�$�!�"OV�P#ƃ�BQ��XA��'7���A"O�[e�ZS�XI�"̓�Jl���"Of�;3B�]�4,�t�ͅN;�%� "O����ωڲ���K4����"OT ��Ɲ�H��=Y�ѵMu�}9"O�� ��7���$�=`x��i�"OL��$	Z��t���2vt�z�"OD�t�������ܴ:�T���"O��x�b^2w��m[�(�/� ];%"O��5(��v"~��H�	���"Oj�:�j�^�
5s�G�8s�����"Ov ��Ǆm�d��UG	�^��ɠB"O4��'�Ʉ��PL�`R�8�"Or�h�+��Ga;� [�l���"O�5� %S;:�qQ!K�v��`u"O�ux����p*F�h�
7\di��"OV���M���f\�x�"m�5"O^x p�C8��h�C�%!�Z<@&"O`a���܆v��l�Uc�s�0 �"O��2h�Q��L��X��!;�"O�͘��S�|k��sFo���X�"OXp��.C�Ű�[1o�,�\Q�v"O8p��R#�D�B�_2�,m�"O��Ȁ��&f����/\	$4V"OJ�h�-��d���Վ9f�z�"O���Ɩm����&;�r�X"O�mb���J,@�F �I�6�%D�,��������@L!�Z���"D�غ� z�.�k@�L�*l���� D��j�oc~���nc ��4D��H4g�2 6���
��q�	r�0D���%Q�7�j�A����X�L�C.D������dlP�c��5-�<2�(D�l�cC��R �a�ꎃj��m;��'D�x ���.Q�K����s9D���������TRp�V=|0�s�5D�c7�)�A�`LL�괮5D�T�d��yG�	�E)ľB`���3D��3ӎ�``)30�@���$�-D�p�c�M42��WG��e�9 ��-D�� J��)J�p��9 �	 �L툡"O���vΙ�vIf �ecV�P��i1�"O��b���c���1��[�"P<��2"O�u�*Ԋz���qL��$"O�- �A	!{u���1�K�u@�0�"OXy*��E�e��!4�G� �*OB�:�*ġi6��  ������'�Bi:��ʄ,,ʤ(���,w=�Y��'� u8��[ B�i�G�`Ր�'���!'��TXR�A'l�ȝ�'V���e�E�ly#g����Р�'֤�NMl��D�? �l��'x���c���8s�C�f�`����'��� ��N3mpXb�a �V�\�*
�'�Q�$�%cz�����T:T���
�'��(����>8��k�� RZ�)0�'X��,Ĕ��TS$E"HS��Z�'$��:0g:h�����D�n<��'�~��dAc�-*�,e��8R�'`�	ٗ?Xn�`��(`5� �'L)�̀IBmBĄ�T}l,y�'8DMz�E@?>p!�X4�b
�'Hlx��S�p���B����Aj|��'Q�uI�	�;1����B2C���'�����Q80�{*ܪh� }��'��@)VK���|�B
��x\���'[.m�v��x[���w(1m�Rx`
�'2 �;rĮN�$�x�΋.)�i�	�' ���g Sq�(�U�ۿ)-ҁc
�'Ӳ�ꑭչ �PS�c�&��UC
�'�֜��H���&`!7����'�Pu�)	E�9q�&K
Ȕ%H�'N��f��;,]���C�J&5�^9��'u��3�Ɛ~Z� �σ�4=B��
�'�*���aޓ:P�9��+��$e�A�'����	�;��as����K�'�<��fJ_�i���lK+���S�'3
$cQk�X.��XB��J��E�ȓN��y��K���ةЧOF2*��&5��P�A>$���Q��Olx��r� �r��%�~	�b� O�긅ȓj(�S���n�+j+�0})v"O�urW��z�(��'�(kr��{�"O�x���D.��� ��P![2�k�"Ox-�ɟ�|^�9�G`ۦM��M�g"O��� �U��DQ��4(�^���"O Xp�-Z�H[�e�E�ʇ0(M��"OD!Q ��.��Q�#�p�Ƭ�s"O��cD�E�Pj��P�ȑL���f"O�ґ)Z${�:�z�j��U��!�"O��j&�V�R��x�K48vQ�""OR��F��3cԈa�ℊ%c�	�s"O�rfl�N *���*4Fٚ�"O���U�Ua�	Hd%]�<���Y�"O�a�,ӌ(s�)2&EG?p��s"O��PF�É?�"$�#kô#&$ܛ�"Of ��n�,b�АhQ�[
����$�=%j�X7�W3�e�B��d��'*��P �W�azN	i��͓_�8�'�b���*�6⺵�E�O�CyT`�'LJTAFᑞWͰٗK��*��	�'��5耍Z�˰9"�j�9��q�	�'/�Y2Qa�m�,%7e4sp8��L�p|�
�6r�[Ĉ����ȓd_�I������ K�@'Sn��S�? R�K�MU�{�*�cP�3Hވ8A�"OLl�"F�B6��S�]�D�"O�uc�I�����Ӓ�@�CH�;�"O�r��(������ow��J�"O����a�M
d�S`���,��"Ot�áOܽ(�J}��f���� u"O.\"�N�?�R�	,2�:�+�"O4zA`ͭ;єh"7���S7�@(�"Ox��Go��ˮx�!��1��h3"Ovճ�E ��~eۤ�=�a��"O�����$bh�P*՘[a�,��"OX�b�]� N �Xj��7+V�"Of�Q@��!*����jF=x���"O��8��ʋ?��B��X�Y"Be"OԌ	Wϋ�J�����	M&W�i�"Oz��܌@(a��M/CqX8��"Of�z6��,�(��/�,�V���"O��P,��]����-��l!��"O�"�� �z�@;Z� 	�"O~���A��)�L�9�J}�"OZ@�p)�Z�B!胂�
8�@q2"O���Ƨ5���z�"�<l�Dp�"O8�8%&K�I��-�T�&H���"O���A��,��	�g�ԘN�bɹ "O�� ��0r܉zr��(uܶhIQ"O��ib�5$l��a��`˾=ɧ"O���N_�&,z�q`.��}�$쫴"O���P��,��#`�&�Z|[B"O�@��M��0^��AA*j����"O�4��jP�i0@��9h��As"O*4���P7VWE'�*d>:�"O&QÌ�6eF�p�eؗNind��"O$���
9�|�`E$٫h�x	��"O1;��P
�4�q���$�"O$��1hөK���1J�;��Q�"OPi�n�
Z�Ͳ�&��$eb�ѳ"OF�0��i�15fQ)#F�TR""O2�����2
4�x$�ݾvH��C"O�"�#. i��B2J���|Y�"O����� )w���c��95jR j�"O(���L�-}@@��н}K�`)�"O��k��ԕE�Q���=n�mi�"O���ԃR~����*��1P��"O�C���:.�xT[��,􅉃"O��p#a��y+f���o�i%N�h�"Opa�C.ATLvAW���M@U�w"O\Y��@�#�h�qpÕ�mZ�(%"O&�����Rq$O�"j��DN�y2(̈n�t�2 �7�	
���>�yR�V�n�j�B'"��z� �9�"OV�YsC2e�Y�bT�� ��A"OR= _!1�a�gP��Vqy"O���q(���v,CG[�w��!��"Oԙ���Qc�L��f9Z��pu"Ol��q`��xS��i҅߾v��$�"O�<@"OΕ&�.��T�Kd	z��u"O��9�C_au�a��Պi���*�"O깠&֮7�|u`�ǣ@��"O|�I�E�T) �D	G=Ұ���"O�0w���|@tsը�9�z$"O�聪�G����
�7�Q
�"O��QwT�;�rp�R �)75�M�s"O���4����â��I��]a"O�iXX��!�|^�1���!�� ��BA�8(B��eM:Ljh��"O�u S��?b�e�B�ѳ:��|ɶ"O�p9�޺I�n������:5��"O�y��˞�B�ʀ�����֝�"Of��c�z8�9�A�"a�-��"OY
��KK<��!)�9��S6"O\!F�$q��A�WGwŲ<@�"Of��d�٭� ���#đT� І"OQ��^%��A� L9(�n`�"O�Ԫ��������� �u(��sE"O�t�#j/lQS��\?V��`"O�z��6t*2���Qը$��"O(�B���fr�+��&8 ԘR�"O.0I�#׮Q@��a�"�?qI��"OĀ���_�	� 1�b^56U���"O\iѢ��+^X�{��h��)6"Ovq�h�9�M07NY��Z�hQ"O2���#$(O (����s���Q"OR�����ln�!Bf��(a�>e��"O(x��.ş�:�d�޽;��9�"O��x��<��1pBB%n���:�"O`c!�Rx&��6�	u�R�
E"O�`���B�8��9�Q���#�r� �"OT�i�.�<!.`��H>A.�tѧ"O�!s��)��5(�I�:�8�җ"O��@@�=�D��Sc��!��9j�"O�13䥓~� L���A�ZD�u"O�!����� ���k�.W7'2���7"O���O�}>LHe��%a0ΰ��"O`)z�E�E�l�I.��|xAe"O~,d�"/&`���%S5\5�'"O�zE/U,�5zp*�|=��I�"O ��bMө;4j�4�$� "O�))��[..�88�bI�27N�y�"ORY����d;J��R���33B5{g"O$��QF���^�{�Œ�=	�t"ON�p��c¸�y���Lzv�У"O�耓��p�2M�T+H"[u���"O4���\/]iĐ�`;0c8�(�"O�d�u���rrm�ff;rPd��"O��9��ѩt��=	��I�ZM,m"O������0�p�U�
�b�#�"O��J����kΘ�At��̴� "O0����ۄ �*��b@a0�IQ"O���b��^�|T��΢L���"O�Q��JQ�F��AD�͹i$zŐ1"Oz�c
Ǘk�NX�Pm��s�1��"O!��V'7e6�j`�?[4�T�E"O���ħ�0��EqH���"O(������I��a�mС}E<�Y"O�D� (ϺNg�@[F�&C��ڵ"O^k%��G��aũ�e����"O:q��B�+-ɀ��_L�n�T"O�Ȣ�B:C�d���Q�Q�h��"O�JÌV�(@(dP��јG�~M��"Ov���ʏ7ZFl3���2a�t9�"O����Rۜ�����26^�Ad"O�\֨�2Z�6 ����EOeCU"Ob�9d�D	mN0� ���!~!Txl$D��	F�2�F�;�h��uwF!�'&'D��£G�u6�p�w	��c�(���%0D���̀�qd���$�RuP�)D��BFL1H:V0P��	(�B��6D��Z���&s܂E*`h�`tB20D�� �)+��Bv�Z(��(� ��"O44���4������} �8Ӕ"O�|�$�.��[��۲*q�]��"O�<���̸X�`��ͣSiԹ �"O��:Q��A?a�D��6kȼ̹�"O��A���X��	�O#�$��"O� c��%�,��d�|8�3�"O¥�g��t��	�''~2a�"O��$iй�U#2h��xm���"O�!��W�� љmM=�B�a�"OR��[;�mj�jϵ9�nl��"O�๓���Cغ����9��II�"O�t�&��[J����Nx���R"O����fі���O��٘a"O*�y� �#����	kb�Z�"O>�S��ǌ!�8�+u�;t�	H�"O�Dc��ŏv�:�A?/�Y��"O�{��H�\��m��N�6MT��"OP�� ,��(H b͘�:5
%"OZ���5=��xa�N�2�\b�"O��
��2.2�љ֏֠P�p(r�"O�U`5�_�g�8� I�t���Q�"ON(�� �/u6�ҥ����q��"O�ͩԎۨBfR<��`ԎQ�NH9�"O@��F������"E.a�����"Olpr�N�^gb�c��3ݾ,x�"O�a�A���tɢ�a��{�
�s5"OB��E�N�&�>�����j/����"O�YhT*�f,���G�6@��"O�	�I9k�����f�?(���"OH4�RG�%�@g� 7hDm�T"O,�G��_���:�
.�� �"O@�����{BE���AǺъA"O$2�əS���f�b�xw"O�;1���O!�}I� _�iJ�"Op,kQ ��1�z��Y�LH$x�"Oj pÌDc�l�� ܩ>���i"O���i����d���M�xo��J�"O��Б�Ծ>���ZBS�k�<��"OPݛ�lV�G`�K�Z�=y�"OJL�e ć�Z1����k�p�"Ob��P,�+�\U�d�j~`(r�"OL����]9r��Iݮ/D��)�"OvyI�o�(�vI��+P�E"Od�(S��;ٌkeєB���"Ot���;r��`�%"*T���"O����`�GWjh���	z�҅��"O(!�g�dS��C�����d"O�`�S"�< l�����P:�"O:�8#��xD���@�]��ȫ"O��37�ޞr��R�G�;��@�5"O�С卄uvh<�3[>�	�"O�͋�BY35��@X5�[�k*2��"O
eha��USeaCW��xz�"O��;Q����cV�gzTA�@��Y�<IŭNo&� Z���$�萨�lM�<a� ���6�D���oF�<�b��9cФk�a\��Yt��J�<9���*V�؁t�^����M	I�<�Cܘ/xJ+��%2��e�ɅD�<����p-@���Ȕ���9��
FܓF���z�K=��j�$f���%�x�ȏj,�:'A�^Ul���D4D����cW�}�,ljbI�"�Y�dD%D�0�f�J:�	��gļ8��X���.D�� j� ���~ܓG��#�~<"�"O6�{��J�M��,2 A
�|���"O|�*��<@�pԱ$nσV��i�E"Oz5BG&ٗob��[A���:���D"O\�3��3yv 4.m.Lr�"O�Yʶ���Z!hC��v���"Oj��'��1� `�qg5�À"Op�$�>?9RppgY�x�1p"OZkd�Ͱ(��E�A�Xs.�#�"O^X B��\r	���ZrP�J�"O��r���_��u�l̈c�ƈ"�"OZ0&Y�-"���VH�%U�p�:�"O���֪7�.u�� ?D)sG"O��!��;AhT��W�/"Z�� "O��
7ٜ=�6H+$�`�� �"ONIA��tg�h����U��)�"O��i�L�(O$E�R/˚f���"O$2���:�Ȉ
�L�?��is"O$peL˒ 6`�`,h²�X@"O*�Hf�³��e��ي7��s�"O�He��CT�e����k�v��S"Oܭ''i$�H��*
< �X�"OP�h
T03)P�:3䅶$��'"O.�8�lȽLU����BJ�p�2l��"OF�;��\��ٔ`�����#�"O��� W�� �C��%;X��r"O��)�׬k�"�)��Ѽu�"�Ӂ"OL �tOY�|����Hԣ�9�0"O,�H�B�!T�<�@'=Q0��"OFmBcԚ|`�GdU=4�X�I�"OJ�#�$�+ġr�"�z�ұ1�"O��# �+-V�J�⚒0�j�`�"O�٠�)���$��o�$�p���"O:4��K0K6��ҥ;׬�0"O<���f�W�.�p���f� ]�"OVii��F�*:�ܻ�\��t�"OJ�ʗ�ɏB� �! �)S|TaQ�"O�Ys%�;J�t-H4����5��"O$�G��EIC������"O�;f�N}��S7��>i��b"ORq�C�U�#~M�QB�==͐ɲ�"O�9�r�.D�4a�g`gҴ��"Oн��m�>��uY��&n ���"O�� �T�=�~t�BaE�9Z�$��"O��L�Tu���`�>6Y���"O�4
*#����ts:���2"O`hjv!G0�s�)��O"�e1"O�h�CG+w_ ��T�ݫf�D"OfI�Q���"�q��	����1"O:���aB u�"%�3��C(��p"O�1��t�&9�6C��*D�Ir"O��Sq����Ѕa@�@*:70�)�"O0��a˃�A=�H��-֘QI�"O�( �>v��8�`B�D"Oh,�FAU�Ncļ��E�
c��c'"O�髖K/;X����]K���"O���w&��J��Z�A�YǨ{�"O��5�V�y�T̻���
����"OD�j��p��p���<=/��""O:�COP��Ƀ �W4�S�"O�@Y&��J�2�x���t��X��"O��A�/�7��x�s@�)�����"O>Dag��"�2�k�iʍ}֞paU"Oƥ���	�e~�m(A��!�z0�3"O� ����gU�U׶0�ԋʉ�z�iG"Ot,C�◘d
,�#����'�,t�e"O*��s�ʊ|(@��Ɏ�z8�"O|t��*> ��FkۄU��,�"O�y���P�<��k�)���xz�"O>��E�b� K���-m��a"O��L&*5�L��鐘4~x��"O�Ӧ��	Q���M�j$ك�"O��YR��>��L�`���Ѫ�"O(u��G҈3�"A{�k��:�N=��"O������ ���Պףx���sD"O���s�^�m�xp���+o��c�"Oh���D��8�b}x���a���"Ol-��RE.�̻3��8d:HsW"O&U���O�-k�R�� S���"O@��Wj�?�LhJ�hP
�l�SC"O��Jųt��Ab���dXW"O6�����.T���XZ�����"O�!ZaD�WF�D�yw��˱"O�:�F�~�1B��̦�+2"OP�Ȁ2a�B�Y��.��s�"Ol!"3@�%F0K	62��Y��M� �yR&
�O¦s�D�0��$Y$����y���/e%L��	ŕ.�I�3��y�.k{T�)�hM�+�<����!�y�G�d0�����/+S�RLZ��y�
)?����N��M��E�b'���y��R�%����mL���aFޭ�y��X�	���h�F��^��҄�y���Ay�p�p�[��~9��V�y"ɘ$^@�P��X��*� M��y����|R�Y�����7�eP�'` �Q��<`�d8���*�^���'D�hHR�֍dMx�s,7�l=��'�,$�T h:��!HCy,@2�'1�}1���=p)|�DoB$�k�'i%���Ӡ�d��%/a��,��'��A�.�fa۠�6em`��'��,�@�����i�n�W��а�'�X*+�5H��d�憛N9v���'��B�mݺ5�v�H�Ǉ6Abԛ�'-�Hѕ��-�H`�킏@3���'f�(:�][�b8�q��"����'7��+5��f̄��	�tb��'�V�č��p5�ِ1���d���h�'2�-��Hګysl��0�N�a����'��,3�	^�*����͑&��
�'vFM�3�4X��Tаj��v�lU�
�'��MР���Q���z�I#o|p�@�'�� ���F=�@���,_!���'62���� �-��U2^I�}�'o��pU̘
 !����ݾZ>���
�'��)I�m�%2�ʄYq T���
��HO��#�N�n�.���!W+�����"OH��r��/v�3�+�7OtL��"O̽���Q�%��0iꏢ Bx�D"O ��>Y�
���II�\����"O�y��h��>�FD`�iKA�l��"O
���)�%P/�m�%%C�iVb!Ja"O�I��Y6n�� �%Nf��"O69Cq��._�<2ɾ�h�c�"Odh�	E�G�v��U�V1,�)�"O��2��
>���' ^$��S�"OF���Pb,q&��`����"O� �5��ۧk-� ��y�j8'"Ou�����E 
Y>>�� �"O�T:o���� �jM��z�Y�"Ojٻ�/Wff�k�j��H٪P"O~�8�D�L)�H['I�*�0�"OР
U1�l�2�ڐn�e��"O���n꒤jw�;+4�r�"O6��&����8��&|'���#"O���5CK�0�xFjB&)�f"O�!�!��{T�E�A�,?hN��S"O�}�JÐp��k�胰kLtT��"O��4O*M�@�:`�@'^:���"O�Q��� E<�e"���Î�F�<A��ZX��
3��8x|�0S�X�<��K�1%α��oNb���i�j�<YA$C
qu�I��RR���*0	�e�<9wo��Vn������t�RDNV�<!��9��Ѻ�/]�u���g�@J�<y�D�(aT�P���
=j�z�"FE�<ك�ئ2'R�
f��	]����& �J�<�1ID�Z.��LQ�m���(�F�<!r�V�>�%��fԇB��R��z�<9�!�q��pu�����aDAy�<a	�q��HX���y#�%W#�u�<YPG��*p�Uv�@�d_�q�R��k�<�!7Z�J^�k�4�s6F�f�<Y�
F�M*��P7���1��a�<�׮N�����/
�δiQB�]�<����:w�9E�������=�䰅�Hʤ� ���W�i�#.�	\f݇�L�Li7j��I�z
@� >NU�ȓ0��A�A�,Z���:�n��2k����E�|��я 6��E��]�����T�C��R�^ �F���e��21x�E��);L�3E�%S�R1�ȓ+<���c��*����7�A��PT��3�h)�bE��cS��4��C2���oтc���l
$v�ȓQ��r'����$p�Q&�h�ȓ]d�B� u�lՋE��S�̈́�8nTSG��!��q�>m�����)������y���3E���1%��\�s��!�ǃ�f���ȓz�9'�N�ұ��֝p�x��C�86kC<Bp.ɫ�B	�[����ȓmj��B5��7����V%g�lm��y7N�X-L�;��\;�B�{�81��[)P���X�AN|�R���	���ȓD�  ��В?p�:!�@�<� |�ȓlB-��Jɠ�yp���!4����ȓ/�`h��M*x�H�'h�;0������e��2�R�g�5�*��ȓ>)���׷&aʐ`5�O��I�ȓ"� �3���b\,��/�1��C8Z�Ȇeļ0���7A[:n}x��.bf\��ؔ`�d�v��9O@�ȓ���;�a��:Q��7=%�q�ȓh逴��#��p���J0�ٺVK*���]u�5���V�&N@��e9S$�0��@�zX��B��n�p���9�P��q������+~M�#�	�Vtj`�ȓ8�~#��B�{>��
�f03	V��ȓY{P8���,i�*U2�ѣ~f���\�d��D�͢B��̂�NƢMf�ć�S�? R�	%�N�t���R�I�zd=�$"O|����4��9K��r��U"O0����+1�j�i��01]��"Oީ�0�[�AwF��c�k�
�d"O%1Gg[�xY�a��*�t �e"OhMX���44��R�i�u�&� �"OhI�bj �=�a6��7�V�Z�"O������^ք4)���/#�؁�"O��Qf���l�v�K�6u`��"OA��4G�}b�e��)p��r"O$�%Iu�*:�.�K� r"O�9�H��D��'ԅ+���C�"O��)�pՔ�3B$��
 �3�y"͗9q���Rpj�c��9k��^��y��Z
2�[�GB.	��ղ�bS��yrǩu	��h`A�%t&H��(�y��Էy#H�A¤L�m�b�{�h���y2儁Ρc�8a�x�������y򁖔�J���脫[>�5����yr��.�8 ��� S�����M0�y��?�h�!�`�]h!�(�y���2I�v�����X�x���h��ym�J��su	U	WHF-�G��y�5Z���!ѥ
�9c��{����y�I
y���F�"����'���y��'AV!�A�5p�) "�>�y��ZF�qx�&�`hh�cW�˳�y��
$�d�jПA$\��Y��y�ː�#�ra���7�61�6�@�yB(W�T�n���)�-]��&���yr%Q��� g� ovjٸDE��yR��3|
 �`O�oX�q�s�
��y��^� 7��;2��PY ��P�t�<�5���h�m� !����R�<�!�@?	y~9)�J�m�R��G��U�<Y��[��m ��A����H�<ː6�����6�4a駫M~�<aE!�X�v��FT�-�t�@Æd�<��e�3�����Z*{���q��w�<I�'OI��yPZ�j�8K�h�}�<FmϐV�$8����r8�"�Me�<���H�ͅJ�0r�؁����ꕇ�j��I��7#wtAG�I����ȓ'0V���@Uj�j����T�w���*��Isɷf�X�c'Hʣp�d0�ȓR��e��A͕n��m�LQ���ȓe�pC�݁AH�#��ڲP�@�ȓ?A�	Qw)͉-�+3	F~�*��.D��X�N^� ��MٱNԆ>"�c$E+D�p���,T��P�սC��	�n*D�L@rI
~H�hD�hN:PR$�-D�t������٠�n[�u>&$XN D��U�X��%�EA�l���XAE$D���4퓈6��	�G�*lհ\Q��5D�<;!S�0��$	 *P9<�����H2D����(��t�`m����G�"`K7h=D��be�
�t��A��M�x���Ad�6D�0Q�܈gB��!/́c"��	3G6D��$k�܂1��M�D���P�?D�(�e@j�����L��,yi��7D���Π@X�A� I:� ��5D�|x�	�F�$�E�0D@��� j/D�Å�� �L�A��B�:!��0A�+D�I�K��q���_0������#D�� ��3�ի5�̂A�qٲX��"Ox�B6�[/G(
p���~�H�q�'�2���Ҁ��MA�*�+nwT�'iX�hfCJw�n���0Ug�h�
�'�����B7[�) dȖ7�И�
�'����mW�1���їP���'�ƴ�D�W�L��Ud� ����<q���`$�q���|���i�~�<���`,6,P�-;�v�ȤO�y�<��N� �h<�B(�%@ ��O�~�<)d�C$<z���pԳ<>|�V{�<�tB�� v(i�f��Nnx���w�<��%5\k&�¦y��� ��w�<��Mɰ0�T���C V! �HCF�t�<��*W8P�r���dt^ 7�u�<�5�x��B#�[�go�z��I{�<I�`V�e?8c3l�n�v�Ȥo�t�<Y�l+ӌ����Լ"4As�H�s�<��7��[�cX򊙘� W�<�5���Q��@;�H� �td0�V�<Q��ҡm�����Q;��ت�I�T�< ���E��(��Ƃ.P�e���D\�<ɱ�ق^����A&�0����U�<��#J�&**��'M՞W����7�Jx�<���D2���q`4a)�Q*� �}�<y�(�wt��(ઁ��d�7��|�<ٶ(=E����ހf�peB��x�<Q����UR½�&��'&�.`�%�q�<y�e �*��@:�)A?�p4�e/�U�<Ä�T�&��r`�&nຕ���\}�<Yu��[+�D�"j˷Qn$}#��b�<��dA�N�$1��6D`D��0ME]�<Y�Kۥ*U�ŋ0#��w�\�<Y���c�bXC�Y��R���Q\�<q�o�3Y�\c��-*�r4I�k�c�<p%�
4����h�Q|M����T�<�ѧ��
ș�ciKt���t/�P�<AFLʰs>�a
�H��g�<��W�<�6엒C���9��$���2�&�{�<YW�ƔyN,M�%fW�I�>��͑C�<�$ ��wl��� K�(|�>LZ4��~�<i�Ø�Tf)Q��R!Jv,|@�#B�<�ubŸ?'�yڠ�I�[��I�fg�<ɳ��U�$��4�TA��c���Y�<)��75��Tqb�Վ���#�[X�<���ΰK~�p�*Ju��z��P�<�T	8ꕱ�l�4MǴ� �NM�<�g���k�@�V%0ER���
N~�<���R�IjD�b!	��N��"�-��<	ǪѨE�d���,��k��$�vmO{�<1R�Ȝh�xlbgoI/\*艹�w�<a㈑p��r�C�a[�=!I�m�<YB�]@ �Qa��Ό��cg�<q�G�ܫ0@�����l^e�<9���rB�ę�&@�P�&��EËW�<�'�~jP���h�i!� �a�n�<	wiI/�I���5c��yp��@�<�B�JQT|��e�u&ԂA�Mx�<9���<و8�ꂜ�(,��}�<I�6O2Ѓw$0}
��p��a�<ѳ��4 ���E�O'ڐ2��Y�<ٰ�N����U3V*�
S�<a�叙E<�pa���@n|��1��O�<��É�$�ɡ�B]�M	2���e�<� �Rъ &�If�"W]�	�"O,9�u� �Qs����vx"OLҥ
�$-4�t@�$��"O�0s���[���&"H���ِ"Oډ�7`۪ �r�۳�_5]j�u"O(I��[=\�2�q�d�
@n�9�"O���fbЁef��P$�d.�-��"OF�x!�[��%�!&
�A��"O�T3��P��<�i�g},@'"OZ�b�CY2=��qf+���a�"O��*�D��

>ty�镳n��YP"O:qR��r,^��h��aܢa��"O�`S�B�/����p'L=�����"Od�I�j¢$���p�=a��}�r"O �B+�-�^I�v�Cn��t��"OV��� O�x���bd	�'
r�C�"O
YVc۝2퀅˕*\�T 8���"Od���n�Ȁ%II?Ar%�w"O�Z���:Kh����V���1"O��� \4M�rE��牻'T!j�"O������$�+1��#4/�"O��� ��bE \���J&�֥�P"O����F&-,|*��3l����"O�Y���Ǳ�p��3A\���|�"O�4�%l!_� ��f@�h�$�6"O`p�f��a8�@�O�dMEQ�"OJ�y4��m���P6�ٷr=v�s�"O
:tl��:$�����+ �qcc"Ot5���L<>��u �����5�V"OD�IWcآ���1SN�)��� �"O �2q#�.�dyB NF�h�S"O�@r��a�a�LeuAx'"O���,�B%�QC��6JH� @"O�@T,�)�0��,��g�`��"O�!� �Ůn�����j�!B����!"O4���X0�pP�̔�+���g"O�L��߭���7�٫Q� �z�"O2�Z��-"̊HY��Ԩ���q�"O�8�R/��	�Yr� �H���3"O8��b/�,T��帒@�\���"O����Q��Ӗ��Yl��*�"O��*&�MH�iX�� �k[�j�"O��L�!4g]�!0|�1C"O^9Ұ�ا[|xiqK�>#&p�Cv"O�4ا�u�$=I��
c��e"O�L��
��5��@pBڴq� �&"O�!��m�T�eʡc���hP!"O��h�o˺�d9�!b�APθ�R"O��(ա֑g���ÀG2E�����"OrtB! (n���Y�@�,z����"O�Sᅐ�,�9����)u����"Oz��f��z<`pãΚ:����"O��ҕ喬S���Ţ�!, ��"O�Dju�B������O���XY�"OfP�]i^䪓nJ	.F���"O����k��
ʪ�#��ط3P!�dW�&�B��6�]������!�$ו(դI�O����p A�;!�d�0K*� X�k͋I-�5I�욾6�!�d�cx���Qm��2+�)�vl�	a�!���h �eP$h%�Zա�5�!�=P�&��F��9��isQ��	�!��	�Vs�-i#	Ҫ`���(�͉0#�!��Xzt�qgT0u�h����^�_!�� Aф��"������1a�Z-`e"Oڽ��DkG �2	C[)��+r"OV1�Po�D��\���M��F"O�3�j�/}���$�F ��}�C"O���ȱh9>P"4���^rH���ȟt��c��]���4�]��e�A�M,P�B��I, #�3��Yi�d�O��CÄ	�F��~�A����<#B�ͪ9	v������"=�v���B7�ؓa�7�*��`
q<䙴	�ẕh��*I�x���$dx�Gx��̱�?A�r.���'��J�ʍه	�>�L��(�w�|Q�����<�|�H<9̗,D͌�K�醄~@:yb�{y2 4�S�DH�0�?�4E���9(Qy"p ��8=8��Q4�nӸY�o�hҊ�D�<�'N�TN<���m T]�+Y 1�.K���1���<��Ҟ'��O�T����_�H�Q@[
O�Ե��MI��M�g-�9e��b"��2����%����h�k��4 `c/ɢb��!T,�.!����F,�?��s����'��s� ���(J��"�,YK�"]�
�ğ���n�IA�'T�	�UZ �d� %� K9��M>A�;O�E����O��ĈʦM�O��7��9H�D�����F3��0R�u-�+Z�<#w�1S�r��?1&�[)Ft�I$N����ZA]r0�f���E���o�b���Ij�Eä!Y���
�/kMD��,�`Pv#܌l���R�'/��~���,X.���8 �-e��'�vy[���?�Řx�^>��'�A��`P�H�B)Z��R$"#L�I����ɥ�?�L�(m4��4��<\]�`�[?�l��ocӂ�O�����l}��&e+���`�;`�����z��X����H%SR�MX�'��哒 �\�S��q�"�{Ѓ�����iS��OB&���	?<�@̸TH?C�x���^��r��b胎SU��qW�G_���0�.�OR6-ӕ���Y�͉�3�2mX��Z�29ش�?�/O�d*�i>	m�pA\�0���;h30iy� � EĂ�?��퓲dd�USKRj��0� �]�D��I�R|:���4��D5C�n���@�O.��y����%\SF0{�'�B���%�Xڀnq���Ifk0V!:�'�M{�i˗!���C�0���01bf�'��!R�F�{�����e���ħIE����P��br#��r�uFzB�S�?i�_��O�&�ٙX
�ߒ!Z�<Ӄ%�W��D!�)�V�I�2^���F��/�h�0�1Y���g����r��aQ'�i�M�K��ix��M�}<��5��:�~b �lo�h��'�i>��W'�G�	��MY�i^m������O<x�21��`��)�Vm�<)��|F{2�Q�
��H�tƘqP\
��M�B�П^����a�z�)��i�rL�A�m >���u�}ӆA�5�'�"��<�SBI|n�a�.T���
���`#^������l����69t�w��:=~�� k\�*�ؒO,t�U���i�ɧ�Ŷ��-��B�z3��҅��6�n�sG�N�h؞����   �   U	    �  #   A(   �pA���d���\�'ll\�0BLz+�lඦ��e�2�<�|:�P��ʌ��,�?x歠t&�6k�u�΄���>1���$4��8(E��Gu���d��h���#��Û��>�MPW�|'+D���s@	�.fJ���Iן�&����ӟ��>�VK�� ���-/��ia�YR��$	M>)V�,=E��;��)_���DK�P�������u�@�4�B�$ɰiH����@t��A#�A��.c��8s�/��\�v����Ѝ 1t�d�Dŉ��!�
of����@�q�Ј����4�az��d�s��#���&M��3Bʓ�o�!����H}{Åw:�� ��'<�O��Ezʟ�[cB[5m `1�8H/z�@u�#�p�(e+���
*��ԥ��[�.�1 �b��j����u�1Od�`�Y-����?�<�!�`��bU��޶p��X=8YYc�L�6�t��EdWWJ��<i����]�I��&�[Q�ձ��!A)!��h��I1���?cZ R�=%�"=�/�x��?���ɕEY*] 1��).�4ks�S���ZdJ��'`f�F���~2�)H�Ë;j �fΚ,iQ� A=��?1�(��M
H���T�С�@��u�<��,^�&ڵx���pRx�Z�A	|�'��y"��9sl����O�8���8�i��yR�� �"eOE�I���)#���?A�W��9��d2��9;k�ZA�z���*�
K�l�{A��0j��f�I!8�c4����o3lr�Q,��t[
���G0����u�[�.�r$
���[$*�&�������R�D��+�MԳU���	@��b�@W�5u�1ZBc�l�@\0ª8�"��S�H�*hy:0�P!8NU"��柌�޴I���'�"�'���'2Y?�rs���Ly�'�?m"��p�9|O�$� �GϓHbN���.��A<�b-�	<U�֍�Ix��u����b�$E{Z�
p�E�h%�S�T�8*b�����%�	�	�8h�i.r��
��-=!򄇶Yj%bV8`�QQ6�3Laz��	i6h.X?%�����D!��W�}+�I5�Es��$�*+%�On9Dzʟ�s2@]� ��I�����$�	1J-�FH��8U�X,~�c>y�R9��pQ���	/8�jN�q���S��2}�Q/w���W�,����	�R�N!�C$RӲ9IY]�b�hJ<�T+����Oܱ�1�
 Xڪ��&lJ��fT�I<a����l��q��U�S�x|���!��J�gBC%]vx���	jX�P�C�JJR8!��G]�z�B�Z�'�iM�1��O -y����p�U#�&lPj�)�)sӌ5#���ʏ|�hAm�C�'&h��v#���0�F9+\0�閍V���Q9`���0��5J �Rw�
�q�i��D�X>ay"�Z�{�K�!mVf0���fp�� �d��t��L<��I�7���rfB�*H�N�a�<�B�� _�P��D�[�*a��`�۟$�'�YA���OHJO"��-�(6�n�2�kD�x���`#�le�}�ܴ%9�p����?�)O�b>i��l̕f�!k�3��p�&�O	�� ��'hXTa�D[�H�
���ÊTj���T'|U�G���9_tH ���q�BD��y�谨â�8G��Iq�F� �	
�ē�?1���'H���r���&�e��Г��y���'T��I��)���0A�]M�
�a3�E<O�1�|�c�O��^�����O�u���<ֿ��.H�k

��5MP�YN��AB�:��Q��"�Xɟ�ӂ&��a��`�C��H�'vh �4hԑ	è?b��	�L��x
0a�!n�:��'RT9���=<���;7T�Y<4D�˓zy����?�M#�i��M�mv:���W+m^�|RC[!Юʓ�?���$� : c����$��+���&��':�#=�O�.�tDN=�P��)L�ڴ��Jh?i,O�3�`��>�p5R�?����MSZwGL��ԩ@U���1��Ȅ��Oz����}�XM��#�73G�	�?%'���v�D+ּ;0�]�h�P��$�)�$��}�����.�ZQ��k�O����Ԅ/$�,��F�;��L<��� �	<��'�ħ_�ٻ�H�e膉�U%���D�=��ð<���VTP ([�`�3V��ac�,&_f#<i2;O^=�Ao��U%�������R��P��XY�HZԦ����!>��0�ʌ#�4��?� �9�b�]�)�q!��ȒUx}��I�h� �'TzLkኙG�Q���k�8�̌�ScŃ@�`� ��
��'J�Zc�)�3�d\#&*z���n],X}5�f#e2.�O���O�u�aM�Oq����5�C��_��Ej��H�L�Z�JJ��x��ʪCV�#$ʙ��T������?��:ObԱ�����>Y5�MAՒ��E=���K�Z_?Qa�i�-x���i o����dB6od��G�ػ!�$N����NX�oh��m�!�D��$�֪=m�h�)��Q�B�ɨ(Š�84瑝.GƬ��l��T���u��$Ţ�	e��?����D`�"=��pG{Zw����p�F�	��
�Zm��n�(k�9�>��e;��	)����MҁOR�Mr1#D�LHkī�"O:� �ӝ��@� (
�|�⠰��'��O�D���H����0�W�s�F���"O��`�L��r����[�L-^q�F�DT���	�� 駄��<G �#Y��=i 
�w�1O� i�O0�0��>����m�v6�� �V�}�6)��L>��##�Q�e�*C��;a�z�<1qO'S�^l� �E�'7�`1 s��hO1��=R��2eA&-�JHi��7D�\�p�/%M�E��o��H%8��@�j�'J���'�fܡ&���Q���e���ڠ�?Y!aM<.�1O�!Z���'�-Qs�@�H"6�+!N��8����J��R�!
��L��H�|�ҍH�	�y�e��Q7���D��2Fm9r�.�O�����;���XwL^�:���"��'>�!��U�.a�a�M6fu�QW�� �>Q��I]̓�"j�-ɢy����5!A�y����v�G�(O���аQ�Uw.��Rn
�U��"f"O�}��@̃g�6rAmO{)�83�"O������]���M
�0yB��¨&4�H��/ �;n�h�G�-��[k1|O:m%�x�s)IP)�`G��j�ͩrc/�	]��u�
��?y�ΟF�8%�7@P:,��\�6�]�]�Rb���c�4��L) �JT��K߈tr��L�l!�$K�NB���ϷUX`8��Q�
baz"��NR2%w"�*{d�"��C�!�ď�]�<��,�)pB(]��O�"j��O4Dzʟ�\ �G�_X��Z�l��4���W8ړ��W�d����d�	�SR���qb�+~w��ʃK�=,�1Ov1tD�Ӹ��r�T5��ͫOv���Jփ7�|���"�\�Y�*̸��SrOڂZdp��<����i�n�f1�P�\5����l��g!�[.�T���O]�!�l�C��V.iD"=y/�T�?1�@E5(��	co]�gh���-������@���'�D���
�	�7/"�*E��O�*Ǆ@S.O���?�eM��� 
&� �ip�+!!�e�<q�f[+(@:�:$�c����HH�'��ybܦt�X]Ї��W�SE X)�y��ї�J��0�L��p�a��?q�Q��ۏ��!�ɓd�������Qu*��t[2�I��M�v�o���O�:�C�܊A��ػ�&��J8	�'�^D��7p��Į�PXb���'�j�fI��f9���TͼI�̕�VO�1J���~(pŨ���+zq1�'�O�	�jE1��
���#�[n���hO�#"N�.ق쉗��
|E��''N���'�4�<�D�n��4Wa
�����O�>z���f��C�	44J�� ��68�nC������;�I� �����̷k�B�ƢA2C.�C䉭Y���� �A+R��AA����ܳ���?187��W�PU�5!A)��c���h�'\�1z*��p\�Q������2#�����{��b�(��oq�ɧ� j���B���	kQ!��'�%�"O~QX���)�\ȣw��9Kf�5z��d7�ŞHu���pk��+DfϔV;Τ�ȓuv�
�	��T`@S}0J)0����|����?9 A���J3yWt�Q�BM0iLb�;�Tc�<d��O�H�p@H�y��x��U�Z����h��v�z�������
!m�	,�)���Oh!��?���<0&�!�H�6�����&f�v��R 0�@Dz�lڸ=��C�	?� �P�Ԙ�v�����q���d�o}B�+ғ��'8q�w$�@nf�26��'BZhl��'.6��Q�b?�w�):�4����'����Vj6D�l�(�@�6Y{ ١~!:�2v'7D��{Ďʨ(l�+1Ձ1\�Z��Ch<�po��,�|�3��"�y"P�T��йO>DّQ�Q1���8@t�d0u%�S��hO���X|b⑐�ViS��e$a��n
��''�M�<I��f�d�<��T��B;4 x�kD�o��C�	`����nݍk=�)�EՍ�b��9�I)+��K��Èaۼ5��ɘ=J��C�	T�9�c�Ա0�D��THV�}ߌ�4���?ŉ�/�b�����oN;-Q�,�pFW�'�b��o'�	�n��	M2h/�}j󡕎%MD��6��
X�.c�1�*Ԋ'Vq��'��a���ȳX���D��&��e�	�'�:<��mס����� ߰��M@�y"�)���6]*H�G��dLަ(:\B�5Z��ꡣ�>VհI�"��,I��Dz2R>)"�i�16c�����R'-����@��?�4��4�1O�嘌��';�P�eeW�!Ҁh�r��+i���IE,̺'�����	��0�WCP+���& !�y�MR�(ylq���R,��Y�e�&�O2��D��C�F샓/O�p��<J�)� �!�RjD�ZU�0�zሷ�mOR��>�#�	a̓�VH@�'�+�-��'a�JH��B���A�(O���+�l�*~*�#c��h(W"O��2e�O�F ��EJ����"O>mk`�.X�fXJ��`�,4�(c��;Zb\��*J�\<H&|O\�'�L�3盌MA<]�Mf���$�"�IJ��u'�:�?Q%�h�0A� ����O�j�B�Pb��+7�7��B o��aS�K�+Yy�I+�a��3�!�d�*|q%x0��_`>T��
Zr�az����%&�|�B	�w@�E�@!n�!򄝹_�0�"4�U� @��)%F�i��O:�Fzʟ��GH��M@Q�s蚉$�~=
P( ������ğ��g�����a^�
� ���1O�T��������^�������v��Z�̉ 6ƚ��X�E�6e,E�J03񁇦�b��<Ɏ��)�Vn�4�"���>�����A!���o4=y�@܀v��@��� � "=�)��u�?Y�2ʐ���P�>�8�ːn����#S�F��'~�G��f!J���E��!�q6l
4;��d�B[0��?��'L3<��s�QDz�����I�<9����%RP��"'u�|j"�DD�'��y�l��l��7o"d�����y��0zh��3���9���r�/��?YpY�0Ҋ�d.�p4�,yU�4Dh DQ�]��	�M۶l�{���O�ܙ0��67f�;w�>�H��':�ȳ�I:0�p��ҳw��E��'a$�rF�(Xaw&�g�Ƶ��O�1h�����0�1�
t��܉�',V�O<�Dܖu�8)�wK�`a�c���3�Ӻ0�B��H�ԍ݇<�����	$�:i�ug<�I 1�1O��������>jt��.E�M��P����y
� 2�3 �O�/�p]r���3LhX��'G�OP��W�D*
i��h�'DLP���"O�UBA#�zؐ2�cEfP���Ds���i�C�n��5J120�[���^�6�=!�dB1O��!�O�k�'�T�S�×GYJd�c�d(8�J�c��L>�עD3{�^8��ٚr�TĨ��U`�<�̍�FG��:a#Ԡ{�� ��C�@��hO1��i��TJ�@Ȅ�3����"O`S��ʹ��qL�/�B��k?�����^�	���##E��a��"ĬL�G)> �	2�5�y� C��?����,g�z<�&�*J�Q����d{�0�	��"��`G�0����HR�>s�͆�Os�9��H�!I��V��'o��|Fx�'�l\�_9G䄴��B�E����'�E� �,7[T�r�!��)#
$��w_�I�HO�c��p�bQ�#+R-� �Tnbupį��޴q��Fy����g��LA���j�L�F�Ҳ�y��0B-�Mऀ��]}����A&�y֛V`<�K!�&Y���0vO@�Ρ�5�4�Hg��P�n�rP�ͦg2�{9����������Zԃu U3$�O�=�;����I�#=�Đ�&�m�1��%�>!�#<��|�В���sa"���=X�ʑ�c�y�"O�X.�>�l���l>A
��� �'I�O@�"�g }H"��K�N�r�k"O蕁���]D�|�RK�0|�f�_p���i�-�zD#P�:N���ÃSd�=i��a.1O��j�O���i��C�,E���W*'�V�s�d��XVI��L>�!Ô0T�M[���*Y�p(�]�<�C�� f��X2�?kg����]̓�hO1��i"���
Dt�ReJ?u	��!�"O�4 �<��@��锩K�<��7���	�m�-M��S`DīKv,Lڱ@�j���I��AA�y"�FC��?����g,$=`w"K��˵�3/�l�	�]�ڔ*wb��M�is""ۮ�!�ȓT�T R�@������(`��Dx��'��L�Be[�P��R�t��(��'��L؂��U�؈F�Ķp�~�{�R�����HO�c�P��%�~uf@@BH�=��� 챟P�4~�z9Fy���һ'2��菾���J�/�y�ݧR��s��]�}�8ͺ�����y�S�S��V�Yw^ɘG.�4F���6Mm�a� ��5�X�m�?�{�o0�D��cS�TL�*�B�%E��O@�=�;q��}��68�Q��$u�t���5�O.��yR�?��K7|���6wP=�E�:B7&цȓa4vqpCU�]�Y�!��	��	Q��,N�b��J�166��i_�o��Ȅ� Ǿ����Ҧ@Lr#I�by��?���)z�+ѵz��Z�dA�??Pi�B"��hO�鲃�Xa�'���S4�F���)�P��؁���:~M���<y#+~�L�>�OT�@�{t�|9P�F��,[�"O�x��� �B`3��P=�.P��/�S�'����n���,`�c��lW� ��n�B��4j�=����DKݏG�����|�T��øcR�h:A�`�0-�G#T��ҊKL��b�p����O�P��B�S���� �?1LI�d�3�
���3��h�6 W�y&���2y�!�$�.�hiu�ͪx�S���!��Ȇ�	1p�jpYЃ�%���sઝ�r��C�It}F\��j�C���2F��X��Z}�I/���'p� �		!j�֘E�y�v���'��6�R�/�Q�b?��@� �dP��!�&��j�g>D���T�F� @� @�ʡc�yň>D�� \�0�?-s� �7��fo�H o>4�xs ���:Yp��͡=���J�>|O �%�8cQ�ڹ6od�A�̏9|psv�*�Ip��u���?I�جV����wFD�=�.�z `NP�4W�c�`��0�)O�Q�D(U�hm�%� �H�J�!�;M��X��b����m+azB�� a<nyj��P�;��r��"m�!�K�ljcL K�Vu��j�+�O�PFzʟ�� p	�'���`m��w���x�<ړ:�����B���㓯)��v��R��y��D�1O��������a�q#�L�c�Bmb�[�Jk|�ȓ,T"@�'̰R�P2���T�Ĕ�<Ɋ��iVW�(�K=s� y�w�l�!��'Xw���G��)l��Bk�>R�"=i-�6��?)iM�	�C3�H�%Xf�:F���MӋ{����bn(�>ap*�(%��Eɖٷ%��]s��i������L}��?�L�;�Km��xr�ى{즹����[0P%�䀺"�B�J��$Kn
��~&�|�C_)v��q���9�̛���7�?��O�=a@����鉮��sġA�!n0ӃlG�u�vB�Ʉ�f9��AJ.U�Z!3gEV�4��I�<�Dn���U�'���6��AǮ��b�ȷ�ϱE��m�B���џ�qR�>���ȶk����'���$1��gL�Z�f�"S@�{\xI"�'4�丗�E�9ü|�l�	��t��LOV��Pʏ� �4��$Jʼ�Q�d?-�Hu6i��tn�0I��'y��j�a3��0H�V�Xx⥀[2�����I���v�L���>�@|��+;�.I�=�d��?(O䬋�'�Ӻ�����?�� �Z�;8��⏉�T��9Ä ��?�)Or����O��Ś9I������n�(�'�|�0-D�HV��
����#˓�D����p-�T�O���H$�腮"s��1�
˓0�����ɟx�'�¸�Р��W����	F���4Ì{b�'7Z�ᢪ�8
��mPu�	H���9��&/�S�$m�(hެ�g/�.]h����� ��'��
k�����%H��'����ix��A����aH�&?�Vd��(�����I֟,r���P�̳�DHH���L<�c��7�4AV�@���a/�$K��8ۥnN��a���UM�ؼL{�S�6����3 ��(�'�5O�k&�'X��S��=qR�N�z��kT$�(�Z�.��C�I�K6�CF䆤�$m	�w���Ezb۟n�B���P�0�~�+��=�r��2*;���� -�d$�(��4��?�TH��)w�K9_pʽ�V��0�z< ��#�(�G�^Rk&.� ��F�F��J�3kQiˇk_�v*��Gx"�'t�%��a.8��5�UMǀ�1�'��k�A�'b�J���@����y����HOc��A&�8���󅏑�*
��un��8:ش �Dy��t�T!�>5����={��P��J��y�'ڑ �!E�}aҦ���y2��.Sk�C�)��5؁��Z����Z�Q�&h�q�x�`�Sb V��{��4�$CX��%K7(�3Έ(Ti���OԢ=��y�L��I�g#���։����s��5G�c��Cr��=\�O~TK7��|�|�@%��;az�;�'`�SI�T2�� �Ƒ�- �p�
ӓ��'�4*u��'( � &P!-�4�3
�'�f\�ЅR�O �ڇB�&,In�i�r�6�S�T�:Bm����]��!�dZ�U'ў`�ta��՘'B�`ϧ9���@E�_�$��S�N��T�)a�yR�D)+����}&� ���$xKD�b�c���i��2D�����3�b!�Ù4sgj�+��#�IK���Oy�A�u���1�)���;}+D=+�'A���0]�u�)HQR���	Y��I4�I��J�%��`��T��� ����N��`�w	�  �    f  4  �  C  �#  �)  +   Ĵ���	����Z�,C�'ll\�0�|r�'~i*���i��� B^(v��8�'���q��+�E��oE��.����qf�a1�r�~X�m��!阽q�D9����m@��~zS�m����q��l;�\0�A�(Qz]@n�$S�A�u�Y�ݲ�$Բ�N@(��@c<qC�"y*���m�8r�ȓ�_�g�v�*�-ݐ� D�#�A� @�Y�G� �Ov 8Wǔ�u'���D#�m�	�"O>	W	NS�q���B�Q8#!�$e¬���A?���+
�>!�#S��ep��_,K��2p��!iG!�$���t�BA`�qh��i%)T3B!�JH1t9�C숊]e�M����'�!�d�`16ik��/Xrڵ����!Dg!�$J7,��r� V
W��X0���$Y!�� V&]Y�Ύ����
�ex!�dC϶i��G�M�������!�ć�C����@��q���ƍڿI�!�$��S"@��UHK|j��ѫ�!�$�<t<�aI�K�[CR��Ӄ�<�!�[�z� ,��X�!�0���'W!�DD�'�)HE�L7)�Ny�5�Q�4�!��u��騣�\�l�t\���-/�!�DN�Ix��K� ����ےV�!���R�hA��6s�b�[�dߣX!�DC!:�(��N�b����ԥ�g�!��2�����Ҫ�br��5�!�䉱[�
u+Ʃ�/皅c�/��Q�!�$RM��0��=l��������!���<!Zě�B��ay�!6R[!�Ě�n�H��%��u<�U���Y�!�d�6�"�I�%�/$�j��5�!�������	X��}�Ԇ,P�!�D�7"p�B �P��AA ��/0�!�D�8�`�§��	]�d�'k�W�!�$)}(9��e�3'�.��U�]B�!�џ�V�a2�@)i�X4�AA�z:!�;ƌ��D��Uܤ�E�O4Ha~�#4",��0�@Q`�`�2ȟ�n�I�M,N�E 4�		3 �8��>lO�q�+�w+�E��K�.�b��	� ����jͪH^�`h�U�al�7�����䎒{[�y!A윊��
G�<yeoY-��4K�x�bU�����<1�f�?k�Dف�.^5y�xhzgkQ֦#}*!��-�N������\�������N�<90.�0�fa�ɇ� ���7���#����o���� K�6��1�̟�t�>YP��@d�(��Ǉ2X���1��x���C�Ԓ*���d�G=��	3΂�H0v1��$ڑl6����H���ȉ� �h�B N�Ii�@L(�R�F|`
�#m~P	��'	M��g�U:�M��X!�ıK Fk
Yhd������ȓe�Us �v㨽�-Q!y�0��g@B h5�����U۸5%rUn:�'_r4 �F�G}N�\ ��� �F��ȓ�f4�U"�]"�0!L�C\}SoN3xe�l$ �"�e����I�X�qj����7�t'Ǌ�r�����I�o`ɉQ��62�h��Ks"i�#�]�D��l""ǂ& ��Ѱ6#���=�!o�]l��C�K��2Hg�'sdm����R9�phsEK2~f�����C�*)� J#o�4���[�<y�!�2�Ե�Q@ǥc�,��H�<�sIU8E�\;-�2@z�z�%��#}J���Y�H��-[?p���W�V�<YGDT�t�0`�)`�,��.�U���@�O�ئ�;h���T�@ϟL�>��IM:��qQ��=�Pu�J���;��`r��Ǣ��&Įxb6�G���3��^lk@�7Fc�4��)�Hș��.o�]�bbG�7\*`E|"S�a���ȩ+��i��C�M�;��B`ȑ�$0`��j�p�ȓn3��[�ϥDS0p��O�V,�̓u�x\K6�9~xk�Ě�Ns�n:�'�r@�c�	[dp�rA�@9'�҉�ȓnĺ��F��e�`���Y���y�D��M$�l�TZ5
��W'��iQe���yXJN�\��w�V���p���j4���F�+� ʘ�b�Q�in����S_��8���ƘE:���/]����
r^j��p)ܺP�a�C��A|">QC�CY[��Z��$L1��r�%�ߦ�ݱ	�8�2F��͈���ۖ["C�		;D(��&� �<���ÐI2���ɿOB���a��),�4Q!qL�7�Ӄ�z�*%�@�ΜqgUVP�C䉯��A��B�.�t�iQ��A7F��Í$(oT7m�>mjP�2��x��O.�I6_����$�,���
7�\pd����r2�;v Q*F�4PU�L���	w��e���c�I�puN)��O؞����*QYj�(�j�|�H��=�^>�UP'.C�0��V閟2��nz�]Q��c7�p�f���j�����k;D��POS�@7�P(�'���)��.D��ADk� q`~��.L�R\�-D��I��2а23.�7.�Nˁ�?D��bv ̼E���xp&&W00�+D��j7-�.|F�s�b[zqD%!��$D��c�Hڋ��S�.�W�$U���$D��f�V�sz�*�*��E�T`�"*(D���@�Q�itQ�����C�v<��#D���p#�
T(���M|M���!D�����$�&�"!&�fF�u���;D�p�g��,��������4HY���8D�D3�b�Mn (�-w�)��*O���h�*0yT9�Vʘ(��H!A"O�$FM^�0|�[��/*ר&"O���ǧ@� �X����\&��Y"Oz�	g�D�	���K��x?8%A"O��{�ѱ%o$Q2AIeH,)jf"O$���k�jt�u:eBȓ���f"O
h �M px���O4*���9s"O8EcEIڲ<��AkR�
�sx\�"O���PD�+HL!��iŠ^qd	�T"O��Qs�Ւik���(ٽEZ�ٙe"OF,@&m�7CBe	��%3W�x�"O��Y�-U�q�h@��ֵ�� 2"O��@bmE�*�J�P� �8���"Od|�� U�T�̅@��Q�-;�� "O�ea7�WΒ�@&V�i��ѳ�yBH��(���xq#��_�\}1��;�yRE�6s"� ٗ��[n��ZF��y�Ό;zs�=agbDM�\����yr�TN���ŊFv�)[E�ݎ�yHK�2�$�P�M��M�4ɒdA.�y`�+h+ɢ�H)L0L�4�0>�������� �\�P��p��a�ΒH�!��T�e��D��낚�hA����R5�O��8�D-ٖ�~B��ޮ,��t� ϟ�qm�T0�ls�<���݀0�D��)>��k�-��
E���dC�I�>�4Z@!Pw��p0i��Px�ȓJ�<Zv-�l��h��ύ*��H� ۃ%W���rg�&��=��J
��k�m�%_���RE�AX��;�nk���gA�nմ³B'�l0�L�ͺ����"=���E�h���4��� u��@�&�(�E�T*9ء��4MB�8D��B�Lv�P��	�}��nL0�yr�ˏH5��{��I0l�`I�ІǺ\W���P�O�Wޞ�2�K�x�ɉ�L>!�% J�XKc'�Y��ի�`�U(<�@;X��ZbNG0-��Z0'сe�\���%P�eft��O�E������:���ct�;v���Pǐ�}�ax��{�ذ1�W�z$����E=����1H��t��҆T?{�|5��OD�Kb�_�����&J�2�4�a��,1S�]�b�h"@˖�;�x���R�'�Ԡ
qM�u@|�1[�,'Pф�更�m��D<�3�+}��HR�F
�9Q�H�EC�9C���3b�D�'��0x��p�fK7�划CQ2u�J\���p�����_'M�U�GZ�h��j�m��t���H58��$�b$ދ��<�`�4u����A�>������Y�x�l��Oz��#A���~W�m2m*� (�4��\X�4C �

d��Ȓ�24��t�Dd9���D��>���8"�(}"�B1=�<�uL��BN�
�$�w�OB��{���qR�mbN�p��
�'R6��D]��Њ���2x�Z&mӫo�Ԥ;������*W������2�}��V�
YRcD�%!r��:|6uk )�WHT�S��^5>}�I�Fr-rщT%}5���� �m��TG�O�:D�3�_�%�a{�B�H�������!h[$C`m�(c�آS�ŵg 8tY�8D�t˰���r�#r�Þ��T���&�	|վ|��%ӆ�>e�,�
U�|��D�ά�'D����٭5y��kBG�-ێ�Y7���X�O�]~�ff���C�9��q��^�(��a�^�s�!�$F�}�Դ!`n�QH�m±���G��v�� ���'O�*�d3i�,:�BN�f 2�U��4�,O�� AƳ�h�q�ƴi/��"O���a�e�NySe�G�?<e��"O.����i�v���"O��R��.B�-�aaπ9���)�"O` *V�-&�1�AϷ�l`R�"OL9���{�bD�kG-3��!�d"Ol��E�24Q��i��D�<\��"O�8"ȅ�Erpdz�%ҧP^���"O��ף�l <���\�RZ�"OL$1$�@�l��#Č�t�.���"O*�˴��PO��x�I��4����U"O
4�6l�S/��ƥF�6���"O H�ˋ��
5��
�&����t"OJ��7�N6"n���	��t�H��r"O�䩧.��MPbk�T��x�F"OhJ���P�Xe�6�ݗbr����"O�K�ɛ�0lNcr�ԫth8�"O|���\K;��`@^�^�6]J�"O���W��#�T�8��ƒO����U"O� �t`Z�q�T��pa@%�>�Z�"O��F�PQ��8"�eH�X�"O���%B!&<���o�&�1f"Ot]��
r����/�P���"O�����:��x��A:��A�"ON�J&��ke��f�eÎ��"O�}�"��*����A��P�İ#"O��`"�N�A^ "2�4b�v̳�"OL�IQaS�k~�AĊP�9��	D"O�AS��(n�7(�nS���D"O���噣G%�,�@d�����9�"O��*��P'
�!�Ꝍ��ڴ"OֱX��4¬XS��*"j�a!�"O���� �'��+�Ĉ>�m3"O�H�%z���pE��#ꢭbt"O&��s�%��A%����X�"O�e(���
�$G-]�0��'"O���哏|�D��saP�|��yk�'8mk�ο8wvQX#�$&��a��:�-��+][@!��ʞ!+O��t�Ȩ�3�[%^����G<�H�ȓK����A�J�pr�`R���:u�"i�ȓL�쀒fø(�Tᛃ,��q��P��8M�0�G�/�}�$k�b��ȓOB�)PfӷC�^��D�2�цȓ}TX��c�����+ A�E��Յ�������]�8���s��)��%�ȓ^�6(cL�63o�pC�h�����g� Xk���JI��Y�-�)�ȓZ�}a��̝c���Va���)�ȓZ�X��2�	;/S��BB�۹ti^��S�? �Y���)Լ4��HV� }��ӱ"Ot��DY`~t{�Y��H98s"O��R&�V~���#��9#J�X@"OZ]	4�F58@�
fn	��"O�Q�D(�%|E0`�ڲq
 ��$"O����*��B�&��qNШ?��"O��c�O�$�f�؇쁄|hQ��"O�Qi�(C�l�x��d,�p�y�"O�-ɒ�O�,����፛U��ݩn҂�~d�PD\X��V��&m�	P���wԨ�%D��jT��)q��-;��f��d�d�"D�xCv�H�\�.�@a&ŹF��C�2��1���)s�lYX��1q�C�J�|�� �9Z�Hi ��4�~C䉜/�(�ccL�Y����a�A��C�	,�.!��JR)L��B�	�j�C�I��V�2g��
x=��hƇ��C��>C퐌��ڭ#�X�`R�1w�C�I<%��Ŋ��¼V����.ݣh̄C�ITEIE�TP�c&	G�Z�B�	?\X����:}k�u�gl�C��C�I�@%	��Db{�)�����bjC�)X���.ɪ��$Z��8C䉍5غHbS#S�����"�V�.kZC�I1~U؁G�1�Q�!�R)6M:C�	*sS�a�M	"̎Y����B��!/���T��vF$\`�a���B�IxQ���V�40E*Pg�0�>B�I�L����x�ܡb��0�C�	�*�B,�F욐zKب��z�B�9h������V����Fľ��B�I�=Cf����C��9P2�B�c��B�	�F;�4P���dR*=� `K1=/�C䉵2�xD�p�H�H�$�A�	ɞM>~B�I:R�\ȣ��V���M���hjB�	�f���K�A��2�T����T-
����)�&[��-��nC(0.!��H��0E�d�׫}��E
P-�!����p�� �&KÌQ��J��!���4�Jd�P��oU���W�?�!��<���xR�FUTH�c�B�g�!򄃭V�f�����E_Xd�����%�!�D�$守�����HG��iE	�!��%���0Ӡ�S�ΐ���5�!��=A�q�J��|��'��'�!�$���d�ZƧ��F�j�3Ѧ�!�!�0PVM;�/�]�v�:G�Ӥh�!�D�;.�R��S�N����Δ8�!�$;W����v@'m���,�&�!�P:Z�~h e�^a ���	�#~h!�Dܯ ��J`�� \≊S�ڬNH!��:+��*�(�46���r�=i�!�D�GW�9����� &K7�!��!`����m��b 4��%�S5�!�@0*h�Se���\|�WoB�{�!�D�ՠX‫.F�<�
�-��!�C ;&a�s(�I��g�V*R�!��[�ʹQQ���M�f��q�Ma�!��V+GĘ)� �I;rT����^b!�Ǌ�XE�ʑXH����5G!�l���P6��34�ܐ�e+�k�!��~t��`>v0F Z�+��H�!�d��#>:!���
 (,��%Ø�!�d�tO`�q0c!z
~Ԣ����Y�!�� v�Z1�Y�r�s"��,B�09h�"O9������8�Ǉ/t���"O��"���3f�x�*Unܡf���"O��[T"�#>ܨ6 �~����"O�|"r"x�b1A#�[�O�f�1�"O�%�ƃ�"���R�j���v���"OPД�R�$!��&��5�> &"Of2��>>`
�y�.��{�,̻T"O>0��
7(��l�A��
��+
�'/�,:-������"�'\Mc�';��J��l���@�*�/2J�i
�'�v4��
�? R4
$�3+c����'��<��i��i�z�y��//he��'ɬ4�E�>kX��Ѵ�\�3���
�'t^̘TBZ���d��;�Z)B�'��=��^�!�� ���,U��	�'V�=���}w�`�2䃮*�b��^�1�E�.`�R%�����a�ȓ>0��ۗb4m8z����y�t��?�����&b	
f��2�`�ȓo�y!���"�d�2FrF⍄ȓPBzdr�[>A��qpB��O�ZY�ȓ1t���Z#n8ar���<�������권N���i*0�[=�l���b��9`E���	~���aF�\�E�ȓb�T)�?C^��#bחyW� ���<�4��Mi��"a�V~��ȓJ��Ij�C�e�p�Ao�� �ȓ+�̣'��"�h���L"�,�ȓ6��}�P���bZ� ��ʪ#�|����4kWo,tٜE��ר�J݅ȓ}��:�G�A`�a��;V(h���B�����K�*I-( �&A4u��%�b�!�a'j�@
&͊`��ȓY.��KS��_Y��Y�Ȕe�*�ȓ.�-Q �?C���CB*D�� �ȓQVj��˘/Ir] ��}P��O3��h0f�	Ey����H��u���'�\	�V��E�l-� ���<�����3�Y��I>C�4|�r��i�N ��	��ԋf��d#�ڦ�]Oj���h����̕(����x�\��ȓ1�B�H[I ��5���\�R)�"O�3C\�&G� �'�27<X��"O@x��/J6�`�z4G��C~�r"O$�U��	�(�;��݆A� ��"O�Hx$H���`�夑��I�"OP��f�Z��Zm8#�/h�[�"Od0���<�(�PĔ�r��:"O�`�J/|�A�Gm\}�D�"O\�j�Q640�U����$�\B"O��#��s� ٢&�;'j[3"O��;vh��np��ą�0ELy�"O<��@���I�T�5���"O<�Л��H��*K�a��}�"O<I��H5u4=���XϒT;�"O(	į
1L���K�^��e"OP�h�D�~h��ɏ�a"�b�"O��r�EW.M�҈2�hO=ON��"O�ɠE�>-�K��.��
�c��y��1��@�IXhl6ǉ��yЁ&�l����3>Y����	�y��T ��}�$�&��2R\��yB հR��5���w����Q��y
� ��4�O�Z��-4�´�q"O0�H��Ƨ��B�7up�"Ol��)\� B���ټq	�b�"OM��戮'fT
c�L�TNTD@"OmR�.]�9$�5�#x[��R�"O�8i�@�I��I���8 �1�"O�IE�ӝ)\F!�����`"O��HP�.m�|2��߽9��)��"O�ݢEf���8&�,Xn} �"O�]J�,I~p,Qa'��KJԬg�<9��3��$�ʱHKL-�vme�<����ʑp��ۯK��Љ|�<i��y�.y�,0Y|y����x�<�c�׉/�>� �	N�<ݾ�X`x�<!�`��`2�ʟm�^4[4N�t�<�"@� ��= ��_��SV	�l�<y��v�*�zcB�쒐��a�<�'�P ^3DQ����\�Jq��@a�<q��^H�+��LdVը���g�<���X�6�2i��U���RG
g�<�D@ʞ?���tA�uV���j�K�<)���^�.�:ǁ's#$��F��K�<��f�TԪ]!RI��d�#�@K�<�u��"���QA� ����ҐL�G�<�6�ف���s���*dƄb�J�i�<gEH��Ñ,Z.8���}�<Ѱ��>G��q�B+��D��YA��S�<	#a�^+���O�k�HY��i�<y�H�l�>�2���-?'������{�<1EkC7Ǹ�s1l� �P�H�iLB�<QV�_$h[��&-���r��x�<�EL�6M�1�����0����q�<�C*��SԤ%�'�$ zq��J�l�<I�	��J
��ԯ��p([eO�<���²q{6���K�
^RE���C�#4sZ�+�H�f�,@�f� ?��C�	�s^(�c��{�T��(�$^ C�I�JN��ARkF��kE1f��B�If�2�r�#�M�(9�^Lz�B��"��e��.�g^*����B��B�	$Vzt�$:�H�j�N;S��B��>j\x!��@ĳo�<͙��y�C䉆&���7�֯�6�c ��<[W�C�ɉ�^�D��!x��j�.�c<XC䉟T�܍hr ������D%�B䉙/����k��v-�����e�C�	���lHG �W�*yK�ō:[��B��48����^�)�Ѓ}F~C�ɅO-�%�#���LF��!cA��=��C�Ƀ{+�ͱ���}b�Yr�ď�c��C䉃	G��õ'� <�tTa�ˍ *rC䉰��( Y��CO�1P]��Ҷ�/D�̱!�������'�E7�=e+D���0gܱ(�\PZ���g��-`(D�$y�F��4-�����:B��e�W 'D��b%>�fu����"8�D]��:D���F�R0��,�,�b�d�l�<aPϘY�a ͢1"��P��M�<�1N#�y��	P�s�48R��BQ�<��"���"��ӥ�g��d�a��r�<����!P!ڌ dJ�
U���/�k�<��EW!6������D�*qzla� Rr�<�!�����c��[��T@�j�<�sk��>����-�>O�)HqeFe�<� R8r0!�r5t@/�"3�,8:�"O
�1#H(�^��#+38| ��"OLԫ��ػgؕ���֭��}{w*O��C��X������f�><��'E��x�cM�#�����M'3��9�
�'�� cE"� �
����[�?��C�'�~!�b�^�T8$a/pi��',��1�G0BL:�$��-Kx��'�(�8�(c21ϓ0$ߤ��'�Đ�u˄3?K0]�B�U���'vΜ���gg��a��C�wX R�'H8L	�R�H�^��pK:&���9�'[�u#�	�=�yj'�A��vT��'�Tp�@ ���   �  B  �  �   S.  �;  �I  W  �d  q  :}  ��  <�  �  ٠  Ϫ  y�  ��  8�  {�  ��  �  ��  �  u�  ��  k�  ��  �  Q �
 � m � �$ f+ '5 �> ^E �M tV �] �c j <m  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf"O�Ya��=!l���Ɔ�b�V��!"O�!)��Y�fx���eE\z0	J�"O>��pg�0Z�2=�C�A�Hy�"Ob\B��;h�`��Ɇ*���S"O�h�T�ÕZ(jܫ� ��+�Ƚa""O�A���I�{"��qReM.v�\�J"O�I��cR�G�Fm+De����(�"Ov�M�{�Ҵ�U���F�T��"O� ��M�g��l�a��8{�Y*7"O�Z��іh��8`�tm�`�"O&ESS��M�,ɠ��b��b$"O,y0GD�!�<�Y#dYF��c"OV�Wc�6�:�3�	�C��:�"O�`y!�������3-�<�"O��!S��3C����ǇZ��\�C"O�V��vA����EE�@�J�yT"OtXa�Ǫ|�t�2&�ۥF<��BC"O�i�w��&dUj��+,1�4�"O���I�tͰ5���߷O�y9p"O��&�(w�̕Z���
P�C�"O1@ŏΞ
f�}KT��}�P�&"O@%����-Zw*�`C�#���O�����wِ;�h04�[�!�� �i�5&֡0U�uy���&�&��t�h�>%?I�U�D��P���v��+��0D������vP� Cu��9M��0H.,}��)��1u� ��7-��0�mJ<qvC�I%o�r����J�1���k�c�5	�dC��#'\!�!�A�Nm��#����!�`C�I�8&b�HU��q�fLr�˜$}�HC�I
/�ֽy���(���K��%a��d����٪ Vč�揗�aN�P��<�!�DU�Ay0����-
SB����Q��F�$%J�(|����i�A0�Ζ�C�	��bP��%���DI��DT�O�7�k��Ip�}��>�4�8i�BD�7@4Qp�	R̓�hO�)���ybF�� =�1�Z�4�$�)�/,fʓX��|���#sG&�����84nY2����'����	�<!0"��2�T�����<*�B��G�@h�<Q ��,������p�Y០�OP�	Z���5/�%��
d˘�+c`�O�-��@�	L ��
 �[�8�!��M��lm�h~]��$?��0/ �q�9Q@�ҖO$t�b#&ғ�hO��J�p��B'�+/T �ao� 6��4�ȓ*p� �ϙ	���a��+4������џ� ��Y��@�BF�`�d:��W,�v��S%%D� ���6,P�ES�hֹ)h:]�ʦ<y� &\�c�����ڭ���9G*�l��	�<q7�Ǚ��]ѥ�.��@���^B�<iWPRN���o=g&�{d}�'�?y��,	0��l�$��y�D>D���q�¯=�����G�04�\q��7D�(��g�Y�0p�*Y�6 	ч͕���x"f��;މcG9d�H���M3�ē�O�#<1c ��L�04�vkQ00<va�qn�E�<Yġ�dWv4#$���veԕ)�*�C�<AP���aX���1���Q��B��hO�O�<�A�o��O�*��u儴<�<���'�Kd�L(WJ.��f�&f��P�'V�u
����x�X�)X�&U��z�'��B$�]�t�@fG��K�^I��'A@�ԉa�Du�u�=�
� �'����cT6Y�pp+ɉ/�t͙�'n�(X����Qjh�"��2-_"A��'-ԩ��`X�5�8�ԫ
)�4��'A��WjGDd���+O���C�'�4z# ݔ'�. KU����\�a�'G����I�3q�`r��� {�Ds�'�i��W�G�T,�Ł��i
�'x|�e�O�}(��yS����'�f�SD�ۙh�HS�I���'U����R����P�j|p�Z�'v�!�O�
uq�lƍ�1e�D��'���u� �8�n��5��0�6���'L��"e�@��Ys��A�'��)�'�@X�D��j���Ç�'�D��'Q.��-W8#�����i�#0��c
�'�ȅ+O�G�x��fR�e�J
�'�����?j^6=A�Y��z`	�'6nU�Q������..�Z�r�'�8��EëD�&� �q28tj�'e�%�W�F�$oZ��A��ipJѐ
�'Vd��P�xQ���@ִkYX�B�'�")��#�a:f}�G3iΪ��
�'T�#�	�9Oˆ�+��
K�s	�'�.�cg��e?T�3����?ƪ��'�@%0�i��2w�9R3�Ź1��DA��� L���E�M~����ǍH4呁"O�5P0���� �ո>;�4[�"Op ��ʠqٶ}s�%
�:L
 be"O�M3�.�/Sny�W���;��{&"O~�AP�Ig�$+1��(/�`���'w"�'6��'�"�'y��'%r�'y�`�6%�3
�-��(,K�1��'LR�'��'&��'��'��'B`l���Fo�2BDD@V(9Q��'d"�'2�':�'Y"�'r�'jJPkaچS�p|�5��%',X<{�'	��'���'7B�'���'&��'^�	�#�9U.�����ZH>����'z��'���'���'#��'B2�'N���`"E4Z��; B��L��D� �'9r�'9�'l��'LB�'���'����S�ΕQ���
�c�,
�r��E�'�'��'���'�B�'���'������I����Hǘ<�5�'�R�'m"�'�b�'���'o��'R1�4�+�	 R$Y�����'T��'V��'s�'��'1��'�2L���Ŷ)S��eE��VbF����'2�'��'�2�'���'jR�'�X3G�O�*F���%�N�jxMK��'���'��'>��'pB�'r2�'�B�p����u:���0&޶�	�'f��'��'2�'cb�'���'hf�J���1�>��A��V���(��'�b�'k��'��'e�jɿ(���'&BU���ܣy�L��Ǭ�>^R���ORh�"�T;t�hʓ���4�dӴ�ZT	Q��	M�`�Ai߃VA@�����I��M��4x�|��?�V�.���w+�R_��i�?A2K�8P���X��Y�m�T�"��&���[�l�D���I�܁�c��T�ZΤL���'�d@B۪a�ao�<	͟J�Z˟�h"��S�,�JׅN/d%ʑ�Q�a�@�d���#1�������P-�=@���E��[�d9�և�?�Tdꉱu�'�<x�F�E�����:gY$�!>=!�`Vn
0;z���O|��+�O�f���G!Gvʓ�y��H��Ԩ���'W����"�&1RA�l�N ��'.�Ip�	�kxs��8�I�92�x��(���b�2oD��ɿJ���������	�(�����d�V�����{��aң��p���k�	��	%�M����riȲ�_l�N��?��K@�4�p��)b�$,�f��6�6��� �<���)�ba� �E��<�(O�(ӶIS�q�@�86b��D0�C�:OB�j�,G'\o�	"�M�G�lD�|�䄘<QD�v�̹8+��ɦ��M�x��N�5�?!�b�5f A]w-���`5O��mZ�4���I1�I��H�	��Vt��J���˟Ԣ�'�&��i�	�����?}d^1' !��5�v�g�ߥz:|�'*Z���.@*1���'OB�O�>��ϟ��#*�?>r����g�� Rd��z}r�'�bQ�~��՘*I���O|�R&��e�"���E%a�
Q�Sц{Q���� %��_-j��$��'���R]�̉�#\���d'+g{�a&�nmH���ԸU�e����?	��?�����dۊyD�Y��OP	D�ͥAy��+�jJ�92U�e=O*�n�ҟ0��)?sY���	˟�v�f�pXqt�Ĭ1挽�F
&P�敓� i�0ul`�h*%o�f��ȘY���.��]7g��MN�
A��m�/x�΍�	ո$R���������?�����R�s�q*���}�vP�l�L� ���`���I֟<����8Mh �S쟈��4�?)���<��L�7N�J��0�	Al@gL��
�ܽ��%� ���ڟ擶.#*���~����'!���1�V1 ��ϽlʚP�i��ڌ���0���-O�1�	
x����V������I��0�ĭ�)�ث��

i$a��-�ݟh��ry"[�Q|Z�c��'�B�'��
�O@"dӀ��fԖX�FGאdI�OD��'W�'j�d��'��!
fh�|��M��^��0�R� ���z�E�i4� oI*�M�����y��h�=�]��+(O\|
�M��k+:T��!�,'��Ag�p{N�u�"��	ߟ���T��ayR�. 
B(��.�0{�Ti�3�X�*��\B �31�剛�M���PA")�'��듀?	7"�&eHB��
\�zN��o��~�,ҊiyjCUCEKZ��ɲ�"�AU��P������yB�H.
�xt��A�B��,� B�-�?Y��'�D/�Sk2�'���O��iqP>y��o�I����%��,�z��O�
��/�������l��d�z�S��)����b�_�= X���1��Ef�?�?��ɤ��2��5�8�@*��u��[�x��5��mҷ"يy���E����1O"��`�?� ��5c�I��?��`�I�=��TMԜ����m�����`��(?:�j���?����?�+O�e
P��>t4���O�DI�h,�`m�!E � s�I�R�~�d�`��	���d�O��05�����cfr�Q�]@��\�T��8�$�s\�I�2�	aw(�ݦ-!�g�r���I;�y��X�K*��M�2D�%�Z.|2@�R!��O&�$�Op��o�I@h��2��O$�$ӈ ��A��Ꞗ�\�Į5<$�d��=/���<y��i��$g��O�D�Nx>u��˪{h����(X@(�H�*<z�� (������@u� A'mT�&E�Z���MY��@�U��i�Ȑ���:����ɟ�t�/�@|�I�����?uj��ռn��T#���;z����2�Y�X�@%�'�d�VE&?��'���O�@l��P��SjَN{d��tf��1��sdCӳ����O��#@P�D�hpT k͟>p��K0u0�`�j

ya �eK�"�� �e� ��D�yI�,��u#�y1U��r��m�@u�'RC�H���B�0�yr�,Q(L_Z؁��?����?	���DL�kjL�%��O�%S��B:��K���l���b�j�O�o���E"0?ѐ^����$K��3R����*��!F♱7���@wPURP��6"Ɣ�a�o�|�q��3V�i|��J_>]�{�? `S�	| Ũa�HX��qT�W�lc�H�a��O����OV�	O�@vR���Ν�u�ʴ� /�PU��3�,M�|����O����,��E%Ľ<���i@C�	�y"�:t�I���ѿ$xmI��Y1t����'��]H	��?�'&tR�_wZ�X��5O&)2�N#E<,����+�hjq�5|,�5J�'���1]�L��EadĠۖ<�?����?� ʟ��Y'� �h��}��霴�?������6-� 
���O����O�����Q�4�(Q#��Ʌ*f`P��#$9%��-��$�Ot����!%�D��:(ҚO�IZ�b�n���X�&A�1��Y���Б�S5_v��C#��<�5H2���4��Q�'+ȝ�ƭ��@�E���V�@>����Ox��F E�t�d�O�)�O��$�<���]EP$x$(D����d
lB��#���?���Ra�6�'rma�O�,�'�RLGS�x�C6o�|��CB6e2+�-q�`[��^+����'�������w*I�jil�	v�q�FW3_�p��qcZ����d�ٟ�j�o94�|��	۟��I�?��s�K{��d��=���:צ�=a�nt�ǐ�bsJ���E$n�	ݟ4�.���D���w�
,���[�yu����I�i͐�1��'҇��~r.]2v�h��O�V0�ո�j�i L#{�ܩ9�@�C����2���@ �i99Ofe�I�<Q��'�l�A�� ����?
@��*7���4��N&�'���'h��36�0��������ʟDr��u6��憘�bZ������
�A??I&]�h�Iӟ*f@����oG��Qj�k
_O4���o�Fn�k�5O�, �����@8TH�7j;��rhR��Q�e(
M�"e4"�←�Jf������?���?�0��ef�<hJ~r��?���i����h��#��!�
��!+�P���4�T��f�ʇ����Ц��I �L�ӼۄY��Ή�C�	!�a��Ο�M�(��*�"�?A�T��^w�ZH4Oܲ� �;�uߴ60��
֡�K��=G	NҶQB��ٕ����Ҩ
�Er`����,���?���M��C��<2g�*.�(pR��܀N{`��'�2����'�2�'���/ ����'��ȁ@��I�2����bFN�
f�>����?qr�O[?q��ޡW�B�(0)��l�&N6����%C�i�C,�,A͢��&�P�<9�]	?�j�d["o]Q�'����Ff�)�K��y�Q/cд�U�]��||�����4�?��?�)O$�X��57۠�D(xn���J�,pX�H����=����������(�Z�,�������u:t��퍰~���b��E�JaS� �'P�V�����?��N`��Yw�vE���]����I���c,`=r@d�Q�tI8�ML�,�|����O����OB�	�|�:���.�'LԲ9Q3L
�,:Lԋ4�O+y~���O���¬�	xe>������q�����	
Kl�cC�6���R��yT���$"��p�w���M8��4���	�(x�M���S�<IQ�� -O�EjȐwϬx�CF�2h�V�S�dx�1U�ay"��O&���Թ?~H�d�O<����B�dm;`��,�h�%�ԫg~�D�OʓO�8���n@��?q��?��\4Z�����T����3��p���w�Z~�(�>����?5�HM?i�"B2:����w�B�Bqf�,]����.؟aS�0�*ԿN�8	�r%�d���韼����']�9�&@�<	%iO1k�l�!���$V����4"���ÐT\B�$�'G�O��'�	����:���(��zC`�9BP�|J��D�<눁�	�lp�4�?-�
�v���ٟĺ1c6A�-�N�V7�+ �I��@��W8t�XA���L�|�I�1�z�����	��ɩ5����QiD/W+�//�	��?a'c��0X&����?9���
aJ��I�n�}��m��?�$�rc���@������?����j�LM���j��L�5i1�g] I�LiH«�W3���O�*D�O#cn����i�����Z�i���.������Jy�F�s'bE�<�J�2iZ��$իwIJ��'4��$T1w ܙ��O�J���*0@`"@�����J�O��$�O��<QB�:���!��?q�R�����(���+RdN?. ����1�'�T��?1�� ER����<� JV��f'�ن���a	8F���I ҚŘsf��n��2��?�!G�O `��8��0��� �rM�w+��O�������?	��-s�
ߖ��'�?��Ӽcp�=FPX�h0�I4k8������?�e�^6uRȓ.O��n��<i��$?�;g�^��!S"���f\�nM��p�,;���1��.m$�!a
�u�gY�(����-ɒ=i_w�J�*&F�9� 2ǧ�	su���&ň Ffxd�'����N�]2e��O����O��i������)Ry�0A/�8qJ��2'�<���|�*O8�D��<S��?��$�D�
�R� �| �$�"� �����O��d�2���\��yyȟ([�� {�*41�� ��A���=����.�nt�d^
)��!��{���б\����9`�	�	�E����U#�.r�J�s��$|xUB���?����?�����9U9~��'�O^Eٷ���%��5�D�SKcB%R���O�n���f7?�X���I����BaV��
M��e�S����.;0�p���v4�QE�o��bgN>��i|ZL�V>1r��G����@ŏF�����]-K4���#R����?!����a,���������&�������$s�tʆ��'�?y���?�VN����'�?�i�2�R��y��t9�m҈�٘�Rل�M��O@�;���[����^���x�) ����<Ƀ�Z:!Jn�����>Bl򱃶�Ī-*�!S�D�O�kF��syr�O�ȧ�Y5s���D�O���=\���jc��N"$�p�(R�-V|��O�ʓU˨ �
�?���?���N�)"h5QjM����:�DՁs�O~rn�>����?1u�w?���P�W�>�S�]���G�Y(y�pT�$i�&����J~ֽ��(��`eJ��२��'�V�P���<y GN�-�ŉ�g�V�+�I��X6�l%�<�1��'��O���'��	&H����D�)wr��Щ���T�Y��j�'�66-�O��3ƞ����O>��;3%Ĺ�.ү:���r�`��SV*���=V��.�5����'�A{��ܺ�bEύ�&�)� ��[���7xP�0!%u�)�'����G�Q킬#�A�O����O��̄du��'*S$hD퍘W�Ш�3���T>ΠrSaݝ%�0R���?)����'��|���/��w3��� "R��t�6��5섐5�'@Ҏ� �~rON8�X�O^��P��B1��Ȍ�j��h2M֞_�jU���B+{7`�Ɍ����5<O�Á�<���'hڰSQ�Cf=�n�+��+��U�^E�a]8v��'���'^��(gL�H��Cy��'*��U�ѕ&�q�4lM^���2�'�$�	�O��'K��O���:���K4hi�ų�:A����P���ɖK^P�!��_?�-�c��|����˟��$hӞs5�� g�(lu^��pgL�Z��'R��'��aJ���;A�O��'4����-0��:��*g[���&���L�2 ��Y���8��'��d��$�&I�i�)!DH�`H��4�Q�B�Aga��|��t�E���۰3+�a��(���A�'G���FF]ĺ#�DG�M@b�� E�6z4T��c�� +%�<��'��T ,�U���'���O�6���@�B�H���ʘ8��c���1�剸	�L$�q
�؟0����d�ӿdY�������EJ�yK�b�xr�
��
�����O��	-�~��R/�j��O�8�k��@>lŔ�@����i�$��,��
��e"���y�(�?T��I�eo8h0)O���+Q�N��qM	/: �b��3]�ȉ��C�*D���Iϟh��ş���Py�_r|8���'�>�Hp�C��*ā&�ɡm�`���'�j6�O��$�����O����O�}���	�4����6 ��g���aak��B�3F�,�y
��|A���My�F�|���w�t!��_�`=�񘷪�#h/�hC��&&�!g�'�B�'��DC�(Rx��y��4ZR4)B�X H�t����~jb�'?�M��l��OT"�}Ӥ�$�"���'U0��7����-*��
4��̲�\��SkW�iݙ�e�身� �?�y��*6Y��׾:>��Ђ޵b�N@��#�ğ�qg���ϟt	����9u^�������	�)�HY��F?� E"�(�+v���I�4�'�� �������'���Oz�\9bH��M���C���8*�ez%!���DI}"�'��ئ�~2��(vg�|�'U�^���,�FB�=���� Bɦ�Y ��A����޴&UK����h��<�rY.����:j��S�$V���q"sn�.Z�<�I3N9F��Q$����i>��Iß��'�$9Ad��;O�0�H��7K��(�!�,6�'�b�k��䔒$��	�����O�lB�̑��\c����)]�Ƥ�O)� G�m4�Sp���`=���p
X{[�MC#��yҫ�%<��,3n�YA��Η�?���'��������'sr�O��Z>Q@Æ׏N!*|��f��Ū��<S���� ���`���m����ı����$�R'j����!��t�s�"�?)�(n|�F~�B�5��`���u�I�(����ב<ǜ8�s�L���2Otu��3�?�Dƒ#<x��1�?Q*��KPƜ��AhJ,	rB*�|xs��X�Bw�����?a��?�,OVĳ��R7D+��$�O,�D����蜝�lI`v@��s����7�	����O�����8�����I	�-{A��>��� #˫*d��0��
��yҌ�0����ҳi�D�/����~ ��:|���Sӎ��5��P����!t��O�������쀔	0?:m'?�������!#+���@�Z]���IG.�V-��{�@ᣎ�韸�	�M���zY���y'$�#a��h�,y%4#3��BnE�bf�#CAr���$� �����a���Ѥ�sK�.��%:T풔&=z����ۈK�����������t*��Ɨmx�����	�?1�F���*���Z��ڷ�x5Х��
9A�p�'�r�9C'�q.��'���O�
��OA>|���[��P�F�p(B#��1� ��?�';��9	��y�3�?Q�r�R��|E��hZ�G���aeʼ[gN8���E�rV��	fX�%�'�Z�P���<���'�l���O���;e��*>�s����$T
��'��'!��'��	�'�`�I��������C9�T�f�,/��Y�tH�ߟ�bݴ�?��@z~Ű>���?�#��$D�'E��P�%X�/�RaS0jɸS��Q�&�I�<�R�6#E�}Ӝt�
�|:��wd�쨖j��?S�M�7$ƍ_����e�0�Xd
��'Z��'}�$��qJ��y'��7c����B-��:A��"Q��'V���$��]�$U���ݴ�?Ga��<��=K�
|�q,�7=���	�)J ���q���!�-��3����$`��1͓NB��K�J�A��`�#��	{*r��m� ٦�	1?5�-�'��dh"�O�Hq����Ox��ڸ6D�	�� �\"-j���e����O ʓsbnje��?���?����ij"%��6��Q&�<Ӥ<1�P�'\�ꓡ?i��7b���'� �#d>I�+R�DXI"�ߵo��*��-�` :&��$N��2�y���Y�bE"�]9Vs���"��s퐎�֥!k��hr1��'�tJ�!a����D�'�BZ��&MO?WP���A.	�`cdQvd�7!��)A&��˟<��+�M��w�X-�'X���?��DL�rz0Y��@!j�:A�����?9�gZ�Q�V�[t�	9T$����N�JW�ͺoZ�&�͓3L�P7,�l�@Ё��Z
w�.$����?)᎓�H�� ����?����`9��I�e�I�F�Fp]�����	}�@(D�]$w�n�d�O����8��9���$�Ȧ�&A�j��S��d���`ʋ84"a��韸H6টH"�$�
l���2�<�;A<�x�q/V���3�G,�v�T/
��y�
۷L�r�ΓV�j��(Ǒ�I�t��SbJ�8#6�ݝ><X���n4�3«Q����	̟��pyr�̤U/2�S�'���'�r,ÓᇤXr(����JHQ��'F�=Q�O�9�'��'p�8;�'�p����-Oj.�$擄O�F��N���N��@VI���չ.��B�@B���*�?�)�!{-�+�g��I�9��áP����K�O~��O��'�7# ������O�Ğf|8Eo��R�҂e�$��dF%�f5s��O�� Ӧ���_��Ӽ���>3p�|�1g�;���Ud�/ 8�R����?����v`�u��<���L9Y�M;
� :��
�M�(���\���Z�.(�I�?a5�ڰj�N�����?������̕Q���S�I\�p8u
W��Y9,OPiX��ӗ$��O�������<��(�#Zd��x7��O��0���ȟD��1x|N�	�[���ә?-��C���H�b�Y�5��#(�72�������P���	>�$+3�'��A�$�<���'ۆ)�`����\���g�|1�.Q49*X9��' r�'���'��I�X.-8e��ßh:%HUz\( DX2ls�Ȱ&%l���ٴ�?1��Cc~��>1��?�t*ڃ���3���#p�h�9^Ly�.��`���V#��<�S�ϔ���=z2�"_>���;k�D2��b�� A
��n5���6�T�c��]���?y���7�ֶ���31/A��H��J<6h\�g�X<�?����?I'�C]�u1)O��o�ПXQ�ac���(�&e.xQ��)�b�hC��߁_�����h-�)��K�O��("��֝�c��4Γ ,�%"7�1Q�=�V��(��)V�^{���n���'���$�6:���
��O����O����C�X)�Ǒ�i]ء�aN�O��<��n�B���?����4�B:��-*�킝3?(��W�?/�|��?TQ���	����&&��|�儙Z�	E� `PD��C��v�����,X<w�T����R?y;�d��?(��O�����v�!{Q��1�|�}���L�$�0�!�?�7O��s],����?�'�?�����i�d�� �_et;c!̤_%��3�??�8���O�n��|Jb(e�4�I�����OP�i���3iy�x��ސ]�\�a�O�8C� 9����T&'A��K'�XY�M[ED��y��՛U��`�Sp�Hlt ��?�v�'�:������RJR�'��O���b�Q>Ɂ$�n3l� �%�AKD�p��k/�<�&�ȟ��I˟���1P쀔'��6=�d2�(�&"��=A�j	�HH�$��O"�dؓ��d؏�"�ɟ��� �i݅�#)A57Ռ8�F`AF��1U�>��Γl�H�q��O��#��Dy��Ov��6�O�&�p�dک2��Y��'K53NT�GI�A�"���O6�$�O�R�cK,�?A���?�D�˃C^Y�O��(�n����8�?q�%TA~���>q���?�")F?��o�"�>A�\��mm��A��v]0El�Ьh&�1�B'�/�j�)�^���'�PuJ���*s���IB�L	\������  ;@��Iџ��	���,�_e�ɟ ��럠��A�l$��_�,d����Xٟ�������	�x�޴�?�1MVo~�w�R����ʐT�8���	�Z�L�C5�ң��,�@�'������D��H�~�4�Ƀ���#վ�RȣG��.�����B�����JNMd�,O�@�	�6ȼ0�A�ɟ�I� �SS��أ� ŋ?���@ɊMմ���Rzy�S&g~�гQ�'�B�'��4�����I�~��\�0��	`9������ 5N}��O����O�q��O^ �P�6��)�ANT�/�3��C�+�6��Ĉi�4a��j� J -3!��]�7�����i�+2�H5�p+4BZ6
Pđ�T^h��[�A���'{r�'��X�AF��(d�ɩp�8�	�~��Y��$��W��	��M���p�'��?��R�l�E#E2ȅG
�+D���1,#t�2oD�P.z�ϓak����|�7m�U�$ʧdg����P��B̌aH��.ȕZ�\ŐR�
Gl��'�2�O��E�����w �4ȶ��{SD����ɞIu���'_-v���O�R
qӮ��S�9��$�\�vm�6b�9�|���U�.��3��O���#]�V��O���k��X�8wgd����oކO��0��	A4 	����Nق%�4�$=O�`���<���'��Y��]*]�b�'��\�P`"�\Hr��颋2A��'�	 I}6`*FRӟ<��ߟ��S�j��Y��ƿ7h�i
q�� Ɛ�k�??a�P�$�����{�,���H��F�R�A�X�8��$Ҝs�j�Y�#֊>����!��i��Y�{\��O(HS��sќ�	WW�����=D� �/_Uܬ��%���?�����!0V����?ͧ�?!���򄉧)�����3[kpt"˓:|�< b/N�U*�2��F�'R���O$��'d���d� b$A3LLUi^�Lk��'f�,8�j)yc�tUΔ��yr�ג#&!���I� R�<����Cͼ�[ŁY�&\���Ɵ��i�%b����?����?Y�'=��ؘ(��P2Fʩm��0xHʠ@5`�s�ʈ|�V� �&�O����O���6p\��#ݛ�w��䁧�=Jưs惗>�X�s�':"d̷�~b��+gz��Ok��z3��:�����|��q���-xi��Q�k&;�I�����'��e�rl�<!��'�F	P��	-�yr�mTʔ[��U�ҩ���,�0<q3"3v�8�Q��?Y�>>|Y�p$��6�N�k�$�d=~\���k֕�'?.��?i��gO����/j��'"*D�Q�CB��i���T�gx��IE|$8�bP��a�0�Lh���[��yRkJ|(��vA-=���y�eDq:�	�I�O8���OP�"��:D���<���O�.�-y��8 #�
4�~Š����c6��$�k� L�TA�O���Eئ��	�Tb�Ӽ�`�Ȱ>t){��4���c���Ťd�U�ʅ�?Y�*��M>Y[w�X)�28O�����u�4?nq�G�,s�U����'�>dCpb»���	㟌�dG��`���ӟ��	�?Uԇ���x$�d���ш�3$��'�������I��S"c���R�9�!��5����3��%\����]���	� �,������Y���2T�dE�U�q�R��W��5v��3���Q�&��P�h��)��P*8tB��	U��˓=�	P�� !�W
�8���$M3A	V91�]����'d��'��X�xy�ǟ�+�(p�ɤk+P	��+74���X.L��D�I��M��G`*��'O���?����FE� T)1��u�"�q�*6J��ě�`�N���3O�q�bÑ&�ugj�<����O�6���8��h3F�B��˫6ٺUcVb�F���YT��O����O��iN��d����Ьc�H�9�1\�L��f ��n�d�O���B:#�����:�D�D���q�Ɍ.�>�	Z�Ĝ�g'FrB��Qb�<X}С�5Ʊ�Tч��>�d�4��ɻP*}�ɊpBB�<	���X�? X\KUiW8/ni��IT��Ă���5�y��V�r+�I��?9� �[�Up��?�;��{���q\��c%�s+�<r��?�.O���B�u�Z�D�O����֝�o����dC��6`C%����91�/?q�T���	�D+�H���� N�H��F2� �S!��%jY�%jS��6dj�A�΄<L�RX��(�Js��OV���jJ����X���0/H;B��`# ��+.�j�Q,��?�נ�&��q���?�'�?!����D-w0x��7�H,*w�,)L*��I���)a��D��V�'(6)�O���'H�b��:Հr�/L��g�)WH��S%9JlP��1X���`�'���3�GӺCӌ��\����> �-"�� �Ɖ��M&ڲ�C⟘�Y�����������\�)o2=�O���H"��D�lQ���[x`�Z�ǿOެ5�&\���	�?�0'?r���yGA��\̐,�5ɂ�|��n�\���'�,�h�'D�=�nTw���(t��NU>^��]� �C� m�x�$ֈJ	|�ѡ+~���N2 J?|b˓G=�헁pȉ�r�'��Pe+-e ۲��@�N|He���'���S��z�d�W�Fx�IΟH�I!#3 ��˖]��k�� [�,�I�uF^�;��IʟH�ɱf3��I�;N<4!��(t&���
� �t�tI0�����$�ahhӀ���/�|r H �<!4"�#V���k�W�����-�l`�'�r�'�`2�G�gt�O���'QrA�:K��^;�ruzT�� v��@�qf�Y��Z��ش�?���E~�w.p=�PN ���Iɡe�l:�"C?K���*��'������	 ET뮀�I|�	�z��x���p�s��$\^M�E�����A�gVH�
-O���I�2��]����ܟd�	��8���R�OX<&^!\V��p6l�dyR��D�TSR�'�"�'	��-���	|��A���h�2�҄]�8D8�'|��O���DV�Ⱥ�F,"Ӿ)�������Ժ�b�:9=��C�M��*���+��T���O���m�Iy��Of�KS+Gy�x�V�_�Q��IC�,�(?���#��O��d�O��$�O ʓD��Ysu@(�?a�����"��gW.��C	��?Iv�i������G}��'�"��K����բ��%p��d2IE��B��'wQ��,P�6��"�d��gl�7�H-#�.�'S��'� p#N��� ��+0��0��$N$`ъ'�ߩ#_��'"2�Osbٲp���w��xPU'��8�5�f/Z@�0��'p�'�.�{ӡ����'��7��O�q��>O��@��:��	�+�
<����.[�6q����&\Y����T�l��)?R�	�)F:qqr��Bu����N��b���'�󄀻mM�˓`S���$��z��'�R�'�vY�tɄ�mx�)*զ�+��'��S����DEhd�	Ο��	�?��g]�9U��z���"��w�.+���qo��֟$��u�����6e��R�O�<��Y�G(�@�Ŗ�l���BC�C���}Au�	-0������֟�ؓ��1����6t�(�h�jC���Y0ș  +��	�,�&�i���x�i>��IƟ,�'�\�D�V���b��)I��Pn��x76�	Ƅ�my"!e�H����5��	�����OZ���e�zn��Sc� P8����O11ӠI<�x���T�x �dPF��[w�H� `��<�2�ںp>�p�Sa�����GC��P(�K2V�a��?���?���?� Ɉ-�� ��C�vא ��O�
Q�E0tK�!^����j�O����O���X@8���ON�lz��y���=SZA��NB�T0��͟��	6Y�~���X��"�?	�S���vN���H@�E��7���@
��M��'[�)�t�\џ���/R�����$�g����|��#½b�n_�6��)���<&HI��㟄��֟`�'�TQ���_�^��'��N�7�����;�<W�Y�E�������d@y}��'����f?Y�F�;�ؕ�f��B�� f�n�p��AE��B�,k�/H�t��˧{+^�I?p�ℋ2���)4�ߓt4� b���B�'J�E�!9R�à����' ��';X�1é�,{>T(�e�
�\���t�'��19 �U3 ��I3�M3��P�b��y�$�SN�{ J��5�rA2l6KO.��t��n �I�}2��P�J�V�6���ɣ-2\�ѽ�4@ĩ�r��F� �\m��(��J�hz*O����/9	@pR�#�ʟ0��㟀��r_JHؔ��^�"��I��u���OyB� ��Pu�Y���I�?��0d':A!ܛM� dH�ڵ*�Π�B��h>�Iҟ��ɢ~D�	)zf6Yk�?�8D"� A�X�tȧ-��Z�M��4jÈ��I)2�JA��'�~�HV�<�v�'U&]bC*N`I�1`�)~%��)��(�" u�'82�'�B�'�I�|�vx0�.��hX4j�V��p��`Իb��͉b�i��9�4�?)���s~��>)���?񰨛!��X�s�Z*0��)M.f���8��K�{X`���<qf.S����_�m��V>	C��	�;cj��(���,Y�̅P���"3NZ����?����"�B�����k���^z2 ü��q���Ր�?����?@��(6��|�'�?	��i���$�y�,� ��H*g���v�����"��W���'"�E����?ͧm��AR\w����f1O�  Z���9AK�7r�M��?4ș��ĶaZ^�,k����(ц�ܝ�?���?i�Ħ���۸4���b���0�?!����»Q�	���O\���OL���%s���c�F,dc�܍r�ᔟ���O��D�O�R�O��(�S7��4��.)A0�ǳe��=��r2D=�MG;�|�`�à�y��o�v���3l'��#-O@�gD�A0�� �L��p,����Z��D�犛���m�I�������`y�W�>t��eA8���e��>{��)c����L_�	��M���a�4��'
���?��b֜e�jYB��Nz����Pi*�d�9!f��P�J�P�T5�:O�a�c�H9�u�fՅ5J$��D��iӰ�'C.do���+�?��@�H�2����?��:�	���邬+b0-��(�%j
���V��Y=Z�V�N�S���$�O��㟪$��,�<�W��y� �&}���K�v$���m���O@X����r��:�����u��6&� b+�f�rTe�Um^!G��1O�,�&�Ԇ�?Y���%�I�?����'?�;�J�j�H`a ����[G�2D	���?q���?�-OJ@�NRK&�d�OX��2B��	i '��O�XI�Ġ�28�� '�������O�ĕ�3���	nl8h�J^�p̰�eo\� ��x*U��y ��Z�tIY0�	F���(�� �U�'`x����'&�L�s�.��b���g�6[D�\����l�I,@�I�橄o�S�l�	�<���$h�%�$�G�(��&�������c�,3�N��Iϟ��4�?���R~�w�<4q)�3�$ؓ񇚽l���3�M�<�r��'w��)�`X\E뮃�wK�扝U�=�W��<���]9Un�B�`U�p$8çȆ�g�2�".O<X�I� ��1c��
ӟ<��ß<�S5wR��1IE<7j����֔X0P����hy�%���<*r�'���'a��Kʫ��t�'	fU&���U���z6.uZ���/�>y���?���HB?)�%O7A��'_"��Z7��ki� #g�,J��]�1�_"sL�ys���<��
����U7!��'�f�F+u�T 6-(��|��ĚF����I.r2F���O��D�O��D�<�Gc�az�4���"�|�A�`�;�TI"��ԮS���"�)#���'��\��OH%�'�r�'F�-��9,4k���/��Q
OS�YB꜠Bkj�h�'�@�0�*�ݺoڳ'�|�OY|��_!N�������o��� ɸ&�~��gFʙt�L�d�O������ zV�$�9��Z�i���V+��[�|�B�"�O����O@�3S�	�O^`n�ؠu�o����i�/4"�i�B��HH��m&�I�i�X�K�O���`[��]"#+���:I���?u4:��"KX�}jީ��J��1LN���fH�'���d�j^,�R�g�O����O�(�ڝb��<
���b��^H��'�ɆF2��Tg����������F*N��	?#�4����٭7��� �5?��]����֟�3�����
��ͬN��iܯT8�S���4*�H(���- @ıH���� "6��h`�韎�{�3Or�9p�<���
�
�8��яKH�2X�nól�¬Zg��	���'��O���'��I�1�!sQe��T��<K7�C4�TkSI�(�Ly���|�4�?yw �<a�<h��ӟ��Umқc��̒�CU#Ba�e�ǟ�9&��-����6/M�����,�ڜ�����s)���y�g�>E���F�H?O��x �*[��?���'�>H��B����'$2�O��M��[>�)@
P�$���{P��
?ՆU���_�!8Tr �����I�����hЅ�'#|7=�Ș1���<?B�PH���������OZ��D�Z��DF�l9��
ȟ��sNk��{�#�D��k�F�&��D�K2W�͓��8Iw��O��ZY,�ʓX�R�**D����'Pj4B�*
�^����S|� 	�b�'��'��]����G;���I�����1hz�26�G?���sB^-k���	��!��	���	(9����61Q�$�E�E�E�	�9�S��E����܉s�6|	��: r�HzS_>mp���O�l��ǫV��a6�և~�L���O�'�4����?i��O�d�!M��'�?y��?��)����8"S�F)ʀ����?�`H�!�����?I1�i��"��4ﰡHV�F/�8�i�k�-n��	P �+\������O6�QB�p�֝���5�M���G`�7�Ow��*a�I4��G��Kk�9�i�<�#�'����dA5��'�b�O`�-��b�"f�~(H���*3�������l7�	)pD��alSCy��'��taƗ��D�'�x��U,��r`�c'�p���f��>���?���I?16'��X�F�'U?��+GlA�hT��5㝙QdI���3�M�S��.�y"꙼��1��	k.O�����P�B���LŒ�CdoXy���!ӥN�������	�����Pyb K.�T����'@`�����T�`�z��_�}d5�'46-�OrL���ԃ�O2����l�íO�O=t1p/ź�x�a�cտVء ^	��k{��蕬��?�n��.lz+��x�ݰ/{^��A��]��՚�S�J�6]�7�N.ErI�	�����?����Pe�s��*D��J�.i �9y>*0�R�4��şd�5��=jfݖ'��6��Oy�3O��dɗ1���s4�])e��s L@Z�d�.>��S����$J�r����%R��	WǒDK�&Y`�MbKz����1dm2�$���(�b6y�0�Q�'��'�E���Ȯe2h��M��n�挣!�'8RW�P�Ahӷv����ܟT���?�`���+/>�CC�t�����O,�S��	��,�I:4Gj�	�N��t�5;�D�pB��FT�EK��6 �F�'c0�p-��Chӄ�{�j��iE,%1�d�>~tj�jp�x�e�6x��В�׎J�Dq1�'Ӳ ��2����u�4��D������n�+sն1+��@g-`���d� ��˓~G�f�'a0(�O��'�ɍW��H" ��o\��qGU�Ɍ8]��3��N�P�D� �'�4��eaH޺�s��>)��	�7YR���f�$JT�@��\t��
�$!�'�	 �y�Iϟ(���?�*-Ad�d�p/�t�q���{�"PK7KƋ���p�̨ ��	�S%Ib�S������K7D��g�(=ہ�V��R��w�ˊ�?y��hPI�1oP9��1²��#�u�CL6F����g������(��\@2�P�>O� �	�yr�&�ɣ�?Q���L�� ��e����g��,�ũ��/(
BX���?!��?a*O�A��D� "�P���O���9��H�ǫ�n]���Vh�0����Q�~�I1����O��ęf���>�0U��e[��ɱF��@Y����y�E���ɪ��s�B�,��=�v�'B0�3)�\�0��q�Y��U�Q��i%����ɟ����_�$�`�HE�ٟl�I� 7i	$p�P�X��d���`%FΟ�2U��!A�h�'Ü7M�O̅�%���>i�0g�+���%/�?D�
萃�V;/h�9�I�[K\Ă6�� k���yr
���;>c�	���ɽNÖi�Â�-bY|r�ۀo;�ʓM���!�D�C�'82�'���$T�BV#�r��˧Oޯ.�.ujeW�0�Q�\8S�\��Iݟ��I�?T&h>��ɣV8p1A�<��]��bHZ�p�y�O����Ov�Zv�Oމ�2�R����ؠw-� rt�.�%1&��nY�5�N$d
R�mT���6O�E�QfF�|�֝@��mDb�a��.���j���Z��q�3�31�t��G�:�p�a1��-�80�S"Nn�R$� x��Y
�@���ֹ�3#��SX�WW�1Y4��t�� �Dˁh`�(W�K���Bh u�L�a �o�Z�kv�E�P�LD+�b�P�|�7�Ʒpktd��LG�5n���J�!F?�����H�d���jd�lÌM´�˭D��:$b��j<�C�ЈF
���РU���1.Ŵ5�"���E�9����fR�&����0���s b�E��M�3iJ�<7���F�?��ʠ��$Kכ��J7�y��':DD�����?��g"�~�#�%��4�D��	>fA� h�����O6���O�ʓ#!
Q )�����'��l�v�ݣ7��ى�мoi��n���<C8B��O��dV:X����.M�Hh1�F��jp���(���nZ��`�	ly���*q?�'�?�����ϛc	8GK�	s�fTZ"�}^$}�4�r��������p�|1���l>�1�ߢ#�X,����q��]� �'���	������?m�'ټ�I%oǌ4
���棚:)�n=;�j��%���'䕁��ć/n��'m���ve�&ǰċu��]�h�شVL�ɩ��i�2�'F��O��^�,ΓF���`�)lax(3 ��7���xp�i��@b���4
1�~�d4h�c)�F{�Q4~� l���	�@J� I����!�$�OLu�f�i��pc(I(tb� �cȜ4<mL�2�}"�R�ǘ'8�'��ÍL���;��Ȅ~#҈��#��C�6��O�͂n�Z}b����y"�'�d�������{Ο'#~LYwF�g���'2��z��|b�'g��'�I�#�̼��7#�$5�����7�:�1D�)��ћ��D�Oa���O���'�r��s��h*%e߆:/V}*�`�4'wZq���'*�	ϟ0�I����'��RAן����~�@h��Q(Uplx��ieh�2��'T��J$�~�'�?����1R���E�g�*��Lc�E8����5�Iٟ����ؔ'
��0t	�~��1zz��&�����ABo�d��T�1�i����~�nJ��?���NH� Q�{򨄝X=��R�M�}C���5�R��M���?�+O��pWÓl���'�R�OVbU����>f���GL�FH��҂L��~R����?I�O����h޽����Yrt�cUF3��@��e��˓!T��$�i_��'�OZ��}E��&�ʹl��3@`��|K��� ���?���&9B��R ҇�ħ)攺�I0u���ǥ[�{6ڱlڹ!4m�4�?����?���9�剞
'�)N�i!,��b���a*���;FMlZ�@N����'���<i�X��ಶ�ȵ{ܨ(��M�Q��!�i���'��@�){�"��<�Sӟh�`�}�|��5#�/-�PP�A��/S-0��i���|�%�~��?���?�5c�M�j$H�3pL9 � ��iX�"�6�h�p�Sڟ�B7�2_�5���{fƌR#.�¨Í�'��V���	矄�I[yRɒ Wd��G�<��������=j�.�<!B���`�	:C]6���?ɗ�u'�98��<Y����l�J��)�޴�?K>�������O ݨ�j�?)�E"��,�����V���Cz�|в���O��
$���O��X>=kQCh�D݁�*�?,��9rk̃�V��x��'�I�,�v�Q�\�M�
B�y���!��<o�v	qը΁x7�&;O����'�P�����)D"��'좡k�i� s���Կ	�p�(��i��R�P��(Ms���Oz�I�?�ؔ<�%8W,��R�$�8A������':�!I���yҶ�0����i����d�P�J��� l�p��>�6j�����?����?a�����	�X�)�4*ڼY����̋	!��R�H�O��ɠ'*Be�U�)�O<.3^��U��.=���A��?��/��*K�7�O4���O<�iTyyD��|�2\:�|i����5G h���ї
W�v'Ip�b�'�ɧ�9O.��G�f�P�hڀ�4��g�w�mZǟH�	ƟDÇ�V��@����'>�ѐ�4EpJ��혃
����`����l�'�dө��$�O����OH�Hb�l���B�[�I�Tu�.�ʦq�IqRѰ(OhA	�O|b#����S&N�z� �T'9��1�F�(3�=��4����O��O����O�ʓ`-���gbF���`�`�|F�pAw_%�	�`���$�O4�0�|������Z���͈�0�
��MS�����Ox��<��^5i�O�)�LK��đhR�|��4,2�,P��y���U?��ҟ�O`F�C�4s�t@2�W�4p�p���@�,'� ��yy��'y���Q>y��K7
 �g��=��Ac��4�N�m�<	G��;G��O��'/��%��H5��,xjB�B�D���Q
6�j�.�$�O����I���4�'��\c�Hp0p�r�@��|��[1=z:�I�5e����O���;�?��S���5FC�$9��rbF��cYP�h�0�M�,O`��D��6ɨ~����
�Z�0�@�Ǒ���8w ]�Ɉ�0��ڱ�z�D�O�10V"�O���?�IQ�ܴ9�X��h�ְ�R�\#D��nZR�4zڴ�?1���?1��2L剴h&��F�f](�&ڐW�V�1bR�%P��oZ,J������H�Iry]>�L�\�����Z��˖�N(A����F�i�B�'���L(t2��'�>��ן���ND�=Ť�2�	�'�L���C�<�8��4�?�����D�u��O���Oh�0ъɪ`t�q6�=�T�!��T�!�	����/O�-��O��C�)[��S�U贼�Uǀ+[��p���D+<{�tC�4��D�O ��|�����O��S���]���Ċ6��ر��=2�dyJ���y�b�E?�ҟ��g�? Čx�*(z*��4�߁F9�0p�ip~��On���O��$�<y'sL�	�T�04a��rv�����N'�&J��yB�'㈝y�'��$�'�Re���.!�����>} �� ������'���'�rP���3������Ob�h��2
����ah_�f૱#M�����i����놡��џ�J��r� �i>7MK�N�"�E�.���4��Yʛf�'q�U��c�����O�D��h�:0S�$N�ᵎ�e�h9���A��ļ�Z�D�O��8OD���<��:�,�ҏ4R<N,�u��2E�s�iZ�I����3ڴ�?����?��E��W����c�^�[1�A�GCG�!�Dx���_͟@�I����w��A��v��a,�,d�*�x���!J�����i��x�q�V��O��D�5�'C��)�'��7�ȅo��:�_�tR i��������'@*������'*x��SMԼ���ܞ;ʲ�㓊h�����O��bY��'M�=��'�"�\0�MsG��6E%\�2���L� ��Ԭ�v}�Z��v	>?ͧ�?���?)�m�@ ��qE
�����9���?JΛ�'����2-�>��-��<I�`�8Γ��1,nqA��֗�` �R0���'�h{�'���'�R�'�Y�l6~�4��4,��qɚHh3+��'�"d# \���q���Ʌ?����?���˟��2b:�I�d�kT����C�^�IП���8��b��'�f̢�p>Q�q��u�ՂS�B�pJ0�mӘ}��4O��D��h3�������Ol]8�W�p��A6o�$j$m�&Z�sC!`Ӱ��O6�d�O*�����R?u�i��r�$	G��8����x�(s�~������g�d�)		����O*ոd9O��'��o^����,� J�L)�4�?i�����6m��$>	���?���D�e��%�*sM�<d���~g.�I��R���O��46O��Oք�;j�2� )�)~A2�9���I��dofy"�[ڈ6�Kv�T�'��$�<1f�18 `�G�҇'vLi�&6[8j�	័(#�`�t'�xXp�&�)-_����Cy�<`��a��Va� �d6-�OZ��O~�IGLy"��?�򅎔�p��0��>���"�b��ps���
8I��|2#ڡ��O�&��8��Ph��9o�W	���6��Ob���O� K��Wy2�D�<y�s�Z=o� (i
��G�.2v�૶�(M܊6m-���^�%>�������	�BF����ۜ.xZ�a[�fE�ܴ�?��"�=h�8$t���O�(�u�?�X�8��t��lW��P�{��QY��6-��ԗ'�B�'�B_�`�bD� [k��As'M�X{2 j�T;��-O$d!�'������i�O�D�/Uk����Z�+ʤ�B�j��[%\�;�*���Of���O���2i1�>���م(���	����'�r}����?Q@�h?�S՟��ɜEKX�ɝ�4@j���M�J��:m�����O���O��D�<9P�ͨ`�O�����б?��I� v��Y0�hv�:��]�nZ�$�|���'�����ʈ=8%���ͥZ,�4S#��W����'�B[��Ƀ�[<��'�?I��=<Y�B�C�G��|2a��,k*����W}?��G�ɟ`��8y�"L��b�	��yWb��j���
���6V z�m��M+O�j�/
��Ѱ��|�D�R��'�jL"tX� gL�i")�v�ؠAQ���?�wu��a���ħ*5��N٪'�ըV��3+��l��uȈAݴ�?!���?i�'M��I7J	����1`��%�6��m�V<S 牳k�f�l��iV���J�I�J�b>����Jܦ�B�b�B^��e�H��2ٴ�?���?12��'%剠XL����O�<:�iu)�O�;�&0�&Ϸ"��e�ش��:���ò����'0�'\���AB�U��ҧL9O=8ex�#l�2�D�P�d$�'
*�Γ�?q��P�\c��h�_��aZR#"F��R�O�]3�m�O˓�?q���'%Kz	8 ��5Gԡ�ꆴm�t�������ɯ|����O�I���?u�I̟`q�+%�优𭚖C��=whƐ#�V���Jy��'l��'*�ɕ4���"�O)b�zD�K��t�)�Z�B����z��	��,�#)���i�O��D֝����գ6pZ�� B�D����G��N��'�2�'(bZ����b���ħ��]��!��W�
�ÐQ�{�i��KK0�~��?����j%ϓ��I	s=��P �C2���� B7zz07��O���<��E�jŉO
���5v"��)�:�r�j��!P��ڤ8��	�+��t�T���?��Zw��\)3/ҟ{���Q�Ǟ{��]��4��U!)J�o!����Od���}y�'�5$�n0�#ݯ�$�T�F�M�����y"�S&�?A.O��S��a��jDF=v�l�QdR�7M�����O����O���<	R&
�|2��8K^R�;P�ӄ)0�H�Gݍ�Rņ
|*ưGx��$�'����3�c�^�@�)$GR����r�b�$�O��MT�Q�'ê-��?9�f�����&d�,vԸI�!6�Ę9�,3lO����O��d�$L�D��@b��7����N��$�6mlZ蟜�r�����D �b�'��kȟk��8sx�!��E��t�F��R�Ҥ(��l��Ɵ �	Ty���(V��9�@��>X|��eZ�Tr�]@��<A���؟L���
Y��'�?���y��!WC�<�0���	ZÄ���Z̓�?����?�+O�H;��|�@�*q���Bڤb�BF����##�Ob��K�(h��O �'K ���OV��͍A�� @�,NTE�0]��	��D�Iǟ���l[�(�I�`��o�th�`�5�$���-�P#��ݴ�?A���t?�������?Qk$�;�� :(����K>����Ô{$4�Ӹi���'�7�"�yJ|����:�d@F<$JS� *�J5ZF���v�pd�'M"��'R��!���ݼ��
�:�A#ꕌ5If5���Ħ��	ǟ\I����h�	]y��O��	�yXX��⅁�tTf��'.�bp��՟̓B#l��w-�S�7T�D8��*ҷ#�
	�ek�<0U6�ħ�Hn����՟�����D�/TLD +>r��e��N�i�$�§6k�7��/F9�����$��ʟЉDKl֙���g��aK��M����?��/��@U���a�O~�$ -d]�6Fp���Kr��Zۺ1ҢC�<��'t�	�y"�'62�'E��`4b��@V��pӭߋYa��)1.h�@�R�J��'������?��([Z�\c��yc	�>���rC�*q�� ��<!���?a����Z�@���j0:?����a݃W� ���ly����?	�L���O��'�����rpF̈%∺v���fK�٘'?��'�W�y�a�'#�5:V+�Wr~�j�W,O*��I
r����OP!�O���'_r��������(M��3�ۢ1�jU�P�Z&V�I̟��	П��'_x���H3�IJ�8�T4���t�����#vf����~Ӗ����t���_����'�2PY�}�� %T.�V!��<�}qp.�:�MK���?�,O�thDoMR�ן,��$%�xY�#
W�1z(��i�z\�Ib���ʑn�O�$�0��H�w4��Au�W.:n�Dp������޴��䖋? lZ���I�Ob�	_Ay�ĭjŜ���GS%�P���O�يz���O����o��@�i*�dK�3���'Ș�>�$x���7���"�QL7��O��d�O����`y�HȦ�?1Q����4���W~](�YW��*����Oj�
��O洺j��'��4�ǎnNB	��EH��%��ß���C���2(O�I�'O���3�M��g��#��i�fG5iw���KQ���<����?��)J�(���C�$��W�Z�H,�@X����/I���|O��ioZ�Wqf��0=Aů��a�͘�X*Y��-��B�I+M��?��?9���?A�Z�������
w���#B�U�����it���g��'�Z��O��L����,���r��\��x|H3���&����ǟ���ܟ���@T���*Lޡ��I�� ��]rz��46�I��?9C�`?�ß$��?�1bӆ�R1�ՋNS �S�+��(�U���Co��sq@�� ĒЌ�vD��2㱟�y�%/�;v�(���ϩ](8�!�"O��S0�y��c��'Q7ڄ�`�O�[��HH
.��a��LY�mъϹO��adaЯr�̠Uً
����g"ʺ���b���|�Iw�	t2z��7B��*��)J� !!�%Ť4���ᅝ�()���X��M��DO:�=����0W>�9���R�*)rq����$���K7�����?����?Ye�Z�oY@�q�f2$�P�@aæ]�rE��JP�0�k�Ȗ7s��?#|y
�l��'a�͡6.�5��<�䄁�����P�<�[(»i+�ȣS��O?�dL��\�c�8c8]"�*D�����e�OB��5?%?}&��xGT�
��,8�`�D���FC䉡I��5òe� #|� r슍Z^O8͓d��9Gx���yB�R���y⇨�]qǉ4>r�'
�k�"�3g��'���'����gg�?KLb�fA�żs�`y�1�C+|�,X҅c�O�p���\�4��鎾����V�o��r5$A�M� �P��dC��I�`7��g�]�=4$)�ҟў�ikP,	�V����T�&%z���T����O�7ړ���N�R=C�F��j���[;	#aҢu�܊D.#���1&5Ȅ��77r~"<���<�-Oؚ&�V�g��a�"ܻ�8�X�M]�[���"��On��O��DW�P�ժ���O@�Sl�:���B��~gt�V�?	�$����5��< Te��а=9�Ě
0�����DC`9�ҩ��6�N�C4@�=l��8'�'� p����?tD
5Zl�m d�بW�ڐ����	�hOd�?�`��	G�h#�&O� �V�\�'��"~�GfI1/=(aL��pPz��4)�<	%�	�<�/O�\X"�qk�D�O@�'tm������=8j4��U�p&A���Pu�a[���?�g��5�Qz� �+Y���t��g-1Ĩ�+I�X����B��z�4�Dyr���t0SvO��j�85�1����޷D�j��[�"���)$D�|�<yt�����\��'��l�5�ń9 
1��̎�#�~\͓��?r���'������,
��F}Re2�S�4/-��dкS̮�`4��&;���& �� A�ll��J�O���|Z���?����?Q��� �������Ja����M�]��E;.�"��'�󩌃W3�c����W��AXq�E(z�ZY�gK��p��X�6��"�ZT�6KX�<E���h ���f��+VB-�r�U&I|L�&"��&6M�O\�o��TG��_��Dy�*
�Q�t��5߶�>u��?�-O����ȍP����5��%1�jJP�'������l�P�Ӻk�OU�a �U(K�̨�!Ih�����'���1�$��E�'���'���I<Oh
�
��'V~����'.,��ac��=��I	�'���2�O��F�yw�����&0"l�@�埌�TaH��`���<c��)� �Aa�(N
Q���R;icx!�e�O� �`��Ox��Ѧ��<)����d 158���F�V:Q�$(�O��1Y��l���"�'|�@m �D%a5� I��)�.¿:��6-2��a�	�'�򤆸}�8�J��DZ�cҧC3	��l3ӇF�~2����OV�d�OR���=J��di>qJA^6z����L�w�d1��W=*����ըw�|(C��DN8 0�=����4�����sL�|r���?���r���%2)K~1z�@�<r���R|0�R苲��Rt#.`C�G~�-+�U�� k��D�	�
�J��V}�]�9bd]�<�h_'8�4����?�/���b��O���@\������ΩX����O��X�Z����&*���?�I�=��0�"o��!U|� �#]�d�<�G�[{�O$4�:Pc�wY�`�!j�$I���A� ��7	���%�'aъ���Z&!}JB�ɉD��1���To<j��B�W8yC����'O��l�'�R���!Аp�"��F�_Y�^t��'�N�B��2�'���0'}����쟜�IP��� 7���/1���D&K�"���*�I}��?yD{��Z�O�r  6���A�Ф��iګJ$����)�矰��̔�^>�L�!�	X�vQ(q��)�DX��w�S��?!�g����� o�&^�֝DF�q�<�! �Ȍ(� G;��+�Th���y��U�O�$1OĤtoʥb���R����Zy�M0)�O��^<_}����L�O��d�O��D�xł���9�bhP��F�][t���4���O(Q��'ξ��u��w��Y�ʈg�9[�'����8�h��$}�!�-�/��,��N��Ix���P5�F�w��<����0/�h�0�<�O>8͓L�p�VLz0��ʜ'z��6�K��R�yBJ�	J+�Q��F�P�$Qp�Y�:έ2�)S'l�'`��'O�p�2�0�@S���Yf�de  X��7ęw��I�d��.�p>	��|y��о?O�u��)w�L��,F��p>�r�]�������w�U�@o�r��64r�B�	:�5�M�	�}�p��{��"?�_@�%Y�4,����ǝ/+^�I���b� H���/?o|)�	�L�O��؁%Xn��cV0v9R��1��|S��P�'Z���!)���	#����&��� `��=[�P	@�νp?Q��r4�/��U�v������g�nl�S�[X�Dy�eߞ�?���i��[��I��Ň7�j�p��?�!�Ĝ:P|�8h�׍N7`��J]l�I�HO�ӓmq���$���"ւ^D�'���)��$Γb>p���-�?�����ɚ�`8��$�O���ҳ"_v��,ĿU����;Uw!R1�Ўo�@ CU�>�x�'"d]���E���[�n�H]�p#�
��"~�I�ZI`�6k�1F*��9�	QK~�դZ�4�<E��a�L�!�B.< (���K�K�$ �ȓ\��u�gQ�a]ƹӰ�\%En�$�ћ'u"!���O��<�p�լɝb�����J�Z���O\B���y�����O����Op�(W��s��N�	="z������	�<��.�����
�}�$U|�(�Zw�ЦT
��p��K�~2Mء��>�2 +��d�������7��v?q'�[ޟD��I4֬H�A�Y6r� �B�&D���]�<A��F
@�x����F&@��y�cɨ+$�Dx�'��'�ΠH�JۆN��и��L�H`E:s���2����'XR�'��͟:�P�b#�'E�IH�/��!��O��y��C���	��ª[H�	��(Ķ��'4�0y`�@�L^z���
4
�D���(�����Ο�����Tx�k�Aа-�T�d)/D�@2� ��b�qA���.���5H:�1�?�U��=V����K�r,~�:�$c� HVh#�I*t�)@b�����z���+L��ja@��UWH%j�g��Բp$�Xr�'khMP��ێtF�L����O29B!FY<<�ܺ�H�Y��`��πB��?� �)�@b��M7�
��	>�{����	P�O7�՘t��/-CvQ���*��i��'ܔ����Ǣ'xl]��"ج���Op�Fz��<�9 ��PA�H@"K@N�K�*_]�t�Ku�m���6�
?d#��I�h�O�)���'�B�']�a��6�Є��U�x���Ҥ
oz� ���H��#b��O�T��@�<��N?��'�&=:�j.EcҔ���X�fJ�5[2�߸E��yS���+�Ri�)��`I��^�h�j��ɓn��O'��U�I����'�?	(O� �ձ�S�ꌹ�cצa��"O�H��-�;\>r��`-�l$�@�x�)f���V�+��?��}-j�@Κ�c<P!ٲ��,At���?�����"N	���?����?��Oכ,)�i��<0�V��_�6���B1���� hd��'o�Y)�ʃ�����	58��`�'Z�1EF"�O�� �rc���MӔx�1x!&�OD a�OL��O�Y���	vyr,�:	�<}�X9d�~,��߷��?	�1O�AHƆ�c",�iB
O�3i�UQsD�;5���)|���'�Z��C.�1h�0i1�o̗j�(���):�ຖ�'�R�'Y�X�q�8�g�'%�	�2)�L�1�O|�9��� � ���ӪF����	�9v⠗'Vb���رC���c�Ɯ�	���p�J-�	ԟ�S���i4�5�'?�pè.D��9��߸N�$(d*o�x(ᴤ+�8?-�ϓ�B�����"(\��Gh�$�3�"�	
(�!�3N�ߟ �	F��/��g@�	0so�.,�p�S����(}0�� �V���'�R�XSf�$J�L��)�O�u�sO��4�,��t$D�:���Ӣ�	��b���c��'�n�ңņ��t���y�'`�����h��)a�ҵ#��U�T�� G��IZ�"OT�I�L�8� ��B�˵C�40�%Y�`��T?�B�;?!äS���9�ѣEբq���<�UB�2����?�)��u#V��OZ���O\�Fa�8����N�(i~�`K��[f�|���E<��ua������\Aq[E�~�I3vծ�CȘ#8���gS�N��4�e���̅����;���S��?���[�k9���h�$�x�̝
l�����?��O�O?�R�<�&���}?FU�V�%Zr"�Ձ"D� ���5U?�E;��)&c$�D��<�C>�Y����(
�H��w�^�)�I7>|Pi������9^��q���֟\��ԟ��I�|�0AAd�P���:���_rP�C�oU��sQ訟��@l1�O�+uL�.F�(qwH�R�1P��O��;�':Tᓴ�R"��M���f�z�3�'�e�����=�!͗�9~�( ���U�0��m؟
�'��"aTb��Y��cHT�A����O�t�	cS@�3�	ƿ-���蕬\����-BP���ܷi\�A�L�.N{\��؝��C�a�>(�ak��i��e��u�Fi(��D&'�P�U�υ�,	�ȓ  HI��HQ�<����0�\��>x��R?�hgßS&�!4�I-�ńȓSt5z⣁E�z����&_� ���z�Ys��#-��9��
�&,�~��ȓg�4���,��:v�!��}���85���)7������hB$���
N$P���/A�de�wD��6����0J9����H���GN�9p1fĆȓ=j�A��"�+�J����9BMJԇȓ ��:I(m�:���'ߴ6R����t��hҋQ�F%/c`A�'�\O�<�iQ���X�@�ɹN\�����p�<!�
y�0h)�T�dxȴ����u�<���F�
"fDjbl\�GgʝR�!Nj�<q1�<0�&��gѲYC8$�6��c�<@"O
e\�@R�.
��<Y�Wc�<��b��$�J쨤�
&�N�oUc�<��)�?G���b�	���- �H�T�<�� Ԏ��P2eS0r�
0ض�P�<ц䕕P��D�E�Fu��[�(�I�<�B S���i���,"<�2��E�<i��y}�]IS�A�3h�BC�<1q_&}*r�(s�УE�2=B�C�h�<���_5f�LL�゜�Z�"�Ba�<�����~��ZPꝖ��i ��`�<Iv�0ܜ*�o̹��C�<�P�s�Ik$�ҋ �����{�<�W��q����tG_�`��b�L_�<AC�J9`���2��f�)A��D�<� �
��[/Lm�����8l��"O��b���@P��ƌ?BL�	�C"O^R���@�0�ʓ?A��E"Op�P�B�=H�d|!�aZ�(���)�"O��(F)�O
82F�Q���9"O�$X\����͂�N�d��"O��9wH@PĠY�b�-x��uR"O�y7i�� ��#cԄD�!�"O|}yDn�9s�R��'"@4{荢p"O@��B��=T )E*ӑ\��"Oά!�G� �`d14I@�f!�P�P"OT��عA	��PC��{��
�"O܅ӣ_O	��3�%H�
N�9��"O	���ԧ9Tt@���'���5"OH=�Å�]!�r��f�X�b"O��AM�=+�	q#̾Lx��3"O�Q�U�B;޼�x�=0o�xK&"O(�����?�h��ǜ]P��Is"O���@ćh�@ ��OM�d4��Z�"OR���ս)����GL(eL*\
�"O0����"Q�0+��ߍ+H�t�%"O��smX���Q�2M�
�2�"OB�c���>�:)���WhH�e"O����lP���(�ׂ�"��$�"O�թt�PR���A���Z�"O�Z#���s�X p�Ĳ$�D�㤝>i����aA�z"�*D��sM�
.#�{�eQ-�p?�KX��
�Ɓ��n쳔`�
���p#2D��Є�?g.�!���-^���$�"�E(�3f�SM\	�M^��أ�	
C�>C�	n}�8�%���\��9DĖ%h�|�	-�Ă����
t���b�϶l1~=JU(��0$DB�	4���Ť�mt�eX�[�E)l�'��d�0"Uu�����N���R�I+Y�;���SK'�O������8�ꀢ6��.Ax�� v"	�e��5�	�'���%a��E�HZ�m_�Z�ּ2��DM-[fH���ɌJM���$����<��
��6�!���G�))p�B��Law��(��DH�'�0
�{�����g�)q�\��<-+��P �!��D?E�$,8�*�{$y���~߉'%�h�`% LOrd����/Z컷%O�h�h�"Oi���$sp,�&](��y�"ORy�p	\ !�LJ����RQ"O���a͓:?���hU8X�j���"OR�Qq�3w�ʆ� �r�j���"O:�K�J���R����L=���>A$f�	��=!�8�r=�2���E0�@ʷ
�w���c�����ar �<
4�lƚ)2��y�m:D���u�Zbӆ�A�fq)¬<�[�I���.DygN/�&�v
Xr�!�D�-1��4Ae���<KJ0@dk�v���(ͤ⟢}�Q�h��Hw$��Xy�<qC��%���,�`��b��V��'Q��!�'�pYk���flh4�b�GH"ȱ�'c��q7	�e �bg��F��'������	D�5a���� [�X�	�'�<��QBh��í�,����'�<ȑ&�5�^�S���3g@��'�	R�B��  ��ާf�6��'#�h���"�H"t#�'�"*�'��`c�.c��T'E2�n3�'u�"f�UX����@',�l�H�'��u��C�2o����&\b�;�',���%G�=�Q�' ~@Px��� �9�#�J�NWN���ȃ�*۸�xg"ON鵇ӧ�y��j��e��iU"O�3�O��#!� j���t"Oҕ�5�x�z����.��}#�"O~���Բ2~D C�` ��w"O���闫V�x+�a��0>fXI�"O����Ϙ_�@9 ��
"#F��T"O��A"E��Km�M�t{ı�"OD%�)�7���͘4U@�r�"O����SL�|��3�hI�B�>�yB�<J��I .�	{��y�B�(�y�阤l�Re��%��:e����y�0.��ez�JY�>�@$F)�yҨπ[����n� �&�����yb.�l�J�iP�q�F �`R��y"�M��A��!�{8�#E��(OR��$�]�T,"}r��*h��V�ܒ/�r@�`QC�<��G.4��p ��6jL$lh�&��~��D+-G�ӧ���߬w �1FNB\��y�t�.��D�(H	(r �8 (�yaT"�y����b����J�G���E�J�F�<3cj�&w��P!�� ff�0��{��MwԈt9���*�,�iWRϴ�`�"��*��H�'���G�0/����D�V}k�)��':F\)#0�� �B�{B�iԵ�y�m�k�\!�����h��8�U��y�M��jŻ�^�h��1�fKǗW_��R��G�k�t���(��M�	�z�����'����ƪ9F��)��i�n�Q�#{��c#C;?1�,=��U"^�H�'���K�Z�؂��+p*�㢚�8�h9� �d>#>�Q�Q�Ȑ�aH�:{L`�:Į�G�\��ks��3.�)�IW����3�Z,x!�w4z4H�w�=��ĀU�'�O4-&-)��\��J��Nsf�q�G�2!R�'�f�s�'AH���<
\tlz���;��AXD2u$J�=+�m�ȓm�Ce!_5���F�R�-���RW���c �
}�]�I�DPX�S6�t�w�7M@aR��+CD��Bq8�0��N�?�a{R �X��ؗ'服"��m�(XW�� 3J*��`��O>��N��5�^2��*�u7�r�'	��B�ºS��8!#Iڇo�D���}���"$�O��� U��c���!=����mz��AD�ʱV�Їf�A^����Ԫt+� SR
\\J�1R�E8H�L�H��p����:��O ����D���� �w�.xXU�70�\�(T���������!�$�!w* �A�ˏ6�D����XX��%�������v�����(�K�?��^�M�4��o�x((R��72D�v/Kl؞��S�S�d���X�xF�&N�U��²dF �Xc~2�гEP��B��h��ƊG`[6+����qtf�) �&r�j�R�8t2�Q�N��`���' �i�'Dqs�>?ߚ\(CB���kV���Ԏ�Fw��{S��.΂\���+�	�a05���@�g��(k$#Q�;~!�cK[
�zR�}�d��}��d���%� X�1��J��� �oO)$����S��Zk|p��@)���m@h�¯�4J>
��vJiy
5DDi�	�WB�<1LD�2(�`��c'L��@���DQ�h�.�҆!��Fk;lO��#��R�Phl�eØ�f0���똔/�0)C���)�'��i�"�0`2 ���Op��M%Ht!e�͡aE`�7mF�g~DI:p�Y�k6P�g	���'�T�[kŔY���S��ћ'-�d�H<��Y�Q	�����J�(rAD���$Q!M�`���!i4"Q�S8�O&0bd�@�.�1b��f�̘ulV��l0�R=gJ�jrǜi�I?cZ扫T�6 �,¢i�
�9���^,�P���(22ؒ���c�`���'K��*Bb[�$G��p�D�"*$4k��*��E�&"�z����3�I���]��}�wJ
6t�B"O�9�퉮�H��+׃A;H��b��*T���1�m�>y�*�BA*)���N=S]��ӧ�+��	��~�G��J$P���I��j*P��k �RX�%���%D�R��-:�I�sDd�K�A�Z@3�"?Ỏ�� ':�t"pN�=Ȑ���ν>��O�vo�3bĥ;ā>ʓ]�����Ğ ��Jai	= ��Q �?H����Ɍ�P����|Rɍ��y�^��ٛ#�Z�2��A�ܭ)Ô�SU�}Z^`�Q!C)\�����˃~��ȥ
�,q1�ٹ�̀�ü=&����a�<�fA�*��P�[���(��x �v$�$MtD�!�'|OBL`�LW4]�~j�铀#�R"d�6rW���_��B)�e¶l!sMо}0��>�'�bI��X妅s!']��1��a^"]z�AC�	:N�Ҙ�&��K�H�4'��n=С�D(�+y0`5��,��@�*Y8�	(O]$������;0Q�� vib��&/�%ҕ �q���� �i�=��ꔖ 2��'�48�����J�1�^II�#Q����#"�ٙ*�ZX�u!�-�
!J��NL?9�ʒ�˰>�a�Z�E�H &F�3A�Z	��Z_��dX���dj�Qਔ�ӛ��HJ�N8�I�j��,*a(�6�h|�1/�6�*��$�rh:���4l���С��08tP�ef2e��<�5O؅å�J�=Q��Q�o�i�S 
?Wh*w�b�'jJ0�,ҧq6m���3&��`&�"RH�t�ȓ2w}��)
"]�@��V�	�a0����g^0�(�ßD�\���M"`g|��z*�����C^���I�by�ه����ɣ ��QV̈!U"�l�̐�ȓg
�sp�N�VJ�A̟4 ���ȓ"r�-�Uh�!b�
��_�g���ȓ;̸��iZR��&	��F��9�ȓZ�rq9&̐�X��V�L!�8-�ȓ/��	���2,5&={#қT#�y�ȓ{�* ���((Q�c���ȓn�b�KG�H�]���QHJ�܇ȓ�z�HS ���!���^��܇��L؂�:W�(m�ԏӬt�Ԕ�ȓN�(�clIG���aŒ([����E��)���ڣTꞱjP+Ң��e��E�A�)�,;���Cb�a��܄ȓt4���7�ڑ|wp�9㢁��݇�qs� �6a"\��ڎ5����0sly��D1�6l��ȉ^tT؅�X�X���ώH��E�!|I��T�������qRɫ�mT5%fц�Sa�2@��6���nJ ��*D�Ș��R�l�P�X�Q������'D�, �L���PeJt�ϮFt`mQ�9D����哇(����#H0w�N�a�7D���rfX�!h� �%m�`�(�s��5D�D��M(K>v<r`K���h��7D���q�J3�ƭ���#���I5D�7��:mu�4�Ńz���3D��Hp���n��!��Y+R%����=D�t���X�5Ⱦ�1�+�I�}(��0D� 1kQ�I�V|��OX�k�"�F-D�@���3�D�k@I1?:�E("(0D���W)B4��8;$g�q�
E�1�,D�,�3�� ;sb�G$F�Q��j�	,D�0����R3f�( ��Zv��zܖB��.�xLk�_6{�4�r� yh(B�I�J�̙�E�'�0� ��S)sS�C��#a5T1��C�+q0�17cFRQ�C�	�z�x�Ґ�)Fkӧ�Ċ86�C�Ɍe�� �
w�.a
gj�2T<�C���*iA'�]��#G%G� C�	i��K��1��ǊTC�I�o��H��Μ�|�f�0Z��B��,Jl��0 V9¤�����B�IH��yy���!F[���!�\$E�B䉮��][�,��D%�A�@k�B�	�b�����셠7*&y�AG�G�B�	�6& ���QdxA��&��B�I4.L�(�hS�+��� p��7��C�Ʉ7�\��F�;�| �Ś�B�~C�*Q6J�P�#�5H�^�i��L�5^C�I:10��Վ20nHX��IT�2C䉿L`�����P�`�VD6�T)G(C�d�l{4B��� �4��cu*B�	�_9�����+N������S�B�}�{4@�%��e�C�2p�C�)� ������_���Hҹi�*%1�"OLx� ���+}r�R�M܍=���1D"Or����T�
�
@���8Z~�H��"O6���!lU�@	�4vsJ0T"O�a;�#T�;��v�'4�k�"O��q��Ty$�@�FD���Hc"O�pK
	,X�0�DQ��T͈�"O���SM= R�0%bB;E��A2"O
@&��0g"]rSǜRﾔ�"Or1:�� �(���ц��O�͡V"O�5!��R���Є�)x�� XA"O0v��>���r�dZo.l���"Op=�f��'R,a!���M>���"O�M�,��yV��u>� �"O�T�# �k	u�P� !$���#�"O�����I�,�q�X�C�|ȩs"O��2�+G��U1 V9/�:�""O��&�P�IY3zP�˶A�v�<q�`���h����
�(_��+�l�<ti]y�j$�kƄf\�i��@�<���N� es�O�uF6�ɅM}�<9��/[7 Ђ��@ C���X�w�<�I�K�p��pk�h�|0X���|�<��[�p��Ɋ§X�fP��{�<2�C�,��e�ǎk��c���y�<Iq��h-���%hW�vG�s�<)���
�zz�CV��TW(�p�<1�m]Cc�hR�b���o�<���5>���['Ù�!�*u��	�p�<��D9b����$j��p���u�<	6CE0d������`#H����L�<�� 
�
^������C�L�A �K�<QR�\�t���G��V��2�"�^�<&/�/�䩳#P>V(��jX�<q��Nd���M֣��g�J�<�4�G�{��5�	?�z�� ��G�<��*��f�)rHI/s���U��C����',@l�rے`������n�D]��'AB9�5!E���"�D��u���'[��iЌ�gM8�) MғX�����'�0t!�	3���Q+e�m�'���Iqc�8B�!��8%�"���'�b��׀��
㤌�S�Ή(���'�&�Ks�W�.nx@r�)c�*�J�'�ց��V0��r�#��\t����'�v�5��#j�(�
�`>$��'6(,&IW� Ȅ�ł
@��	�'6��h��['Ğ�P���/_�A		�'-Ҽ�oC/}^�t;EEʂ�6�j�'߮���n�9Ԙd����`���'U���'ҺL$EH@�j��(	�'�̔k!�I0,o���f	ȴͪ�'��ݨ�N/J�Z2H��c�'�JͺwjE�]�Z90�`]�t�Vex�'Q֬����0��}���o�r�J�''X�SI�7J�4
֨D*y	r���'=��VCK ��s =DF��'p�kے6a(�b#�5E.أ�'`	ȇ�N�r��š/&]J�'���" ��Xcf��B�< P*�'�bq���A�.�`�4Ȅ<����'P����ÐA����@.ܲ�,�1�'\�rʑ�d�֬�@oG�Ґ�KN>)�n���hY�l�
( �+���.�y
� �i��d���G$V�G��'�'���
0� ru���J|�f���k8!�$��|h������3+Tu��]�W6!�${�B��>$2���*�!%>@��'�j��UƎ���A\&-D�P�"OvL�S��:%�*T�5�N�$v���"O�`w�5O��Т��8��9#"O4�)�c��!�-:��+���"OL��'�$A)��2&D,��r"O�PA�ؙ���b���y%yF"Oz4�!eƋ������(`G֠j�"O}۶�Y0j��\�� /ᖽ�B"OF��� ��~ Ʊ���_(	$H��O� ���8$��*"�D�_�2eH�g�<QwJR6YC^m�@J ^�4��p�Z^�<!��N�B�l�b�i��^�f=It��Y�<Q�葋s��P ���5O�����}�<yFl4��4YS����M@�C�T�<�@��l�3"�
�pٔ9��
Yv�<adi�D��p��>�t�BN�r�<asK�H�b,�7��+ޞ��An�<iR�L�(:4���b���̻��!D����`���g)�qPb(�R�!D�\z��0���:1c.�2ˀ�=D�|�� 	�Zw1��Y��0���':��t���'^�������?Pqԡru�L��ȓoj�xF��W�j�2!��"���ȓ*�,������\��aN#u���ȓ@���0�>^0�*Q$�t*a��5�<񭊝&j��1�~����ލ�SoGd��W��$[~0ą�~O��ȡ`M�&+�� NM	�D����J�@�/ݏ�\�!�F�	�ȓdl��G�	%�4�g虾BZ�ȓ~!n Җ�]�uB钅�ǔ�f��ȓd]J�#���?9�rSE�Ї�p�}��"��}�ӆr"ԇ�2e�Pakʢx��т3�BH�j���C�,{� ܑtD@�:��A?P��ȓ�.�z�h�a��4��j.g���h^��@�'H��֭/|�:ۀ�a�6E��@ Z�QX,��
2�=!�ċ(W��+A�������IN�Hr�Y�U��I�4��Q $��hޤ3v
0*��싴�B>~80�?����~r3ؚf�H�;GO�%Y��k�I�e�<I��3x����2� �|��V�=�䓻�=I���a(`$jA#
�=�3{�<A� P�T���'HҒ�zH�S�^s�<��;yx�k�EMC}�D���OF����>顃�o}~y�4�R b�e
y�<�藸G���[{7�����|��hO1��z�j[�5�\%��E��v9� "O�9W"��� -���x�Ό��"O����1w�Pd ���� D���gc��T���2��!'m>D�P�P䑷 6��)��94���d���hO�4KP1O>mpDY:;
\�A*s�D���"O���ŉw���� ^;��,	��DP;/��b>m��KY���u2cF]�<�f!�b�8D��������nظeM�qY�o.����ia��R����c#Í>��1f>D���ã��
Ӕ a!��䰹��:D�x��_���M	A�k/|irc�8�Ik؞� a���`�,�N����%�c"O�P�6�{�`��w$_��l�C"Oޱ���]+3] M�D��= ��5��"O�c�^1�V��o�Yn��I"O�q%�T8.E�BdM>R8�"O��{G�ax�0�cg��9�"Ob�(t��P�8���f {�"OJ1�f�J����C�/6ED�8D"O>���j[�[xf0@�A�-{?.%X�"Oia��ǂOk�1�k[474y21"Oιʷʏ�H��a�+L4
'x0�"O�I���A.B	y�D�.|H��"O�$���èP��) � 'Vg�*�"Od�j�̗�+���A�Tf��0S"O����bC6��=QW�(:q�"O�)��H1E��c��)0��r�"O�h��ll3�ݨQ.l0�W"OvA�d�W���;���w�Q�"O�Q�" ��zQ���C�mZhq"O\ 4�W)KF^Pcs�S�6�@�p�"O>���mм1����恜w���r"Ol�P�Afd����@�Ү&�y��R3�2���,
 ,�^=���З�y����%�Ĵ�&fE*n���fn��yBJ�Aq���a��8:`���Q��y��C<Q�Bx�A/_�@�aO��yrF�w,X��!π|/�p�E��y�L#FPAҖb	�p68���!�ym�4v>>4
��Z c�؁֩�yRI�_���qb��V���2��Y��yrO�b�X×�S-N�h�!$-L&�y�^�dƼ��
 AvFD("����y��D1�	��:���Cd+Z6�y��K�
���x&�I;9�8�	��۪�y��O�5 h��sA�35
x�Q�&�y"J��� ��Vc�&�Ҵ�E��y�L��l����E��\6�ŀ���yr��+B��ZF�Ψ��T��y2�g{���FK�<w�je� �͘�y2��wU��8�Eذ@fp񐧂�yR'�6:����1�ʷ-=�ɷ�Ȍ�yb����
ʎTf�-K�DV�y�ߪX9$EC��ùQ�Y�	-�yBW�3j	��5B��a���y�F�8s:�%�_�9��Q#ף�yb��F��j��+�<���F��y�G���V�U~�p �ޚ�y���a,����	I,�2�d��y2��VrT�1f�[�HS���F�-�y2`��N<QY �DI`Nd�6�K#�y2-'O<
�w��k����b^��yR�:@�)h'R�6�"��E	��yҮ�E����)(Z<�#�â�yB��"=i򤑅Q&��(c���yB(��F�}���ӦNh��*��9�y���=Vj�ɓ3���1,���T���y�oK�9c���K]�+��Ġd���yR�ߒx���Ff����s���y��G�4�B���)��3��y"#�3����`#
�-��Ρ�y�jW�*�F�jg.���`�|���PG���d��
&��=`��U94��Ć���)��E�r��Q�'k�.)�p1��X����/�t���A��)h,�]��S�? ��ZJ��d�xҢW�(�"O����Lw�� ��kZ��&d	�"O�@  N�6�܁a�KW�D�b"O
�Q���D�64�k���=�"Oҩa��0ZV�H�oF
�R6"O�Բ %�#A'`�fh�� 2~���"O@�BbL]�<�D�O(K�p"O���TȒ���YH�F�4�q6"O�U����
n�Q�ʋsZ�"O0�L�g��mC����DsR��a"O>���V�wb�yq��o�-�"O����R$s^x�C� �Bh��"OX�����'r�T��c�a*�z�"O�e��	f�h\���vh�"O�R�J�;Y�")�ã�"��}(�"O��C�ԬH�N��`i�.P�6��@"O@H����~u� �3�|	D"O����b�C�6L��8.���"O[���MY`|�BeL�4xD"O���ڛ �|tdS2[���f"O��9󊑯@���Tb��D'�y�OV�_� ����Ң�tr2�:�y¤�=T��%��+������Ǣ�yB�O`2q���Xu4�rW�y���z�`Q��Aܔ\9� !Wn�8�yr�W�@�I���"R�M�����y���\�&�[� \�J3�A����,�yB��-h�M[ŏ��+"�<�&O��yB�M�+� S��T(��P#��y��Ȍ9����K��&��$J3�ybA\�zネ�d+�#o�y�]�O�ʁ��ۙ��$��K��yB%^rcp�)u��!fI��@��y�]-H\Lѱ,��e���\,�y�Mҹ?�^�(T/���- �L��y�E�d��@f�C�{<�pQ�V��y��\�{�Z�j�C˫^�`M�����y�*B*B�� ʓ��f3N,*�m �y�Λ7���2�	�Y�@�b�]8�y�4�d<RЎU�g�T�ѢG��yB�1�>�a"�:X��`j��̷�y��11S�S�f��Qĥ╠Z�yreC&�R��Y�%���!
�0�y2oO0t%��B�o*$��׋�yroZ�.���j��y������Ԍ�yb#�$zY�u#$,ξz����w���yr�V�_e.�"ӭ�s������G��y2���M?��@�AEg�x�#���y"�N�]�VШ7�Xa,�e�:�ybĉ�S.<�[�O��Y���y��4�y��Юk<��PF
M��r�jUʚ�y��4b.� ���c�X�+��y�
Њr����BF[&v��'�K�yңâ^�v���?Ô�٥hJ>�y�-�&H�ĸ�*Jm*8�����yȒ)��`L۪F���K��y�iU!wqH�#��!>�!�P��yb)�1��t0��8 �I����yr�^�kB^�"�N)Q�� U�F�y��6z�t�q��d-�',��y�&��e�F9i�@�P�ļ�����yҠ
�?4��RB w9&����0�y���ir� ze�[/ ��Jr"�:�y��^Φ�X��۰����f��y
� �l�oT�j�B����|��"O��A��˔f�00gI�'����"O��9���4��`�ES�!�>�#�"O֌2�����cS��Z�ȓ�"OЕ�0#��FY�!�1�Г`"O$�f^�y͎��`��~
���"Or��b��?���z��$G�QSV"Oj$Y/H�xwJuR��֜�I�"O�@��ơO��)�e_�;��8"O����B7px�S�<"��Q�c"O��:cԄ�P��u�'
�dH�"O�L��+�-��-yL��!n`LPd"O�ip��ɼm��4�ш&`-�@"O�
���+_�äLN% V�l*�"O����M���(ܲ֡8@'(({G*O� `C��)����(4ZK
�'*��I𠁘U��sV��6*�a	�'$
:��Y�r}�-�UB�4:�PA	�'�~!�C���K��9�'
�aA�'�|1�GʝQ���#M8fP���'��@�$KM�(o8�x�J�VL`y�'�J�ߦ{�)�!a�� -꽐�'�Tڗ�%�`�gEǫ	I+�3D�Pe���^�D�Z� <��!t�#D�ܩ2L۬]L�;�m�+H��!��#D��#��S�v���囦_
��ka� D�2�c.�v��A�=��09"n>D�`	��m@�Qr�<,LJ\B��<D�(c6l�!'(��p.�'�� A7�-D�H:"f�A��à���>��x�*D�s��A���}Ң+�*��9�gD;D�~3�KՠɏX,���U��A�zC�I�e�0�s��q�${C�Ӻ�C䉛"y�t�X*l$p"�nE7`�`C�ɥk��R'a��7�<�J�D�e��?ю���=
:��q���6�:�ka��7z�C�	y�����d���0�qM�
�C�ɲ,�4,k��^>c�h�k��Md;�B�?(����X�rX.��G�L =��B�Ik3dI�DF��f.q*�KP�Y|B䉉M�^a��M�J�Θ�q�L�A~DB��2Ax���Ь�-bd$�X#�[B!�lK��TYnq(g�-�b%��'���"�A/4\A�֏ѻ��	�'�$@�bP�O�@���eT/�/'D�0��-6g+��1i�"4����vN%D�t�0��$]�b�ڇΚ�pC��9�!#D�زD�W/>и`WBX9*1zD)�O=D��j%Û)�j�x�ŗ*'�N�K:�O��BR`=(TIͽV�n��4�rC�I�6j����SF�$��#��[u�C䉅3S�1S�섇-b�X��9=��C�>^�*�(���S&$lr���;��B�ɺ+�r�`�'H"F���q.R?-�C�	���2��j�u�$�۞>8�C�� T|�R�+�Lł���Xu�����6�&;��b��5Q>��Aؼ/ǲB�ɾnr@)3�ꉑ-4�Y�3�S�C�B�ɘH��]y�n*!9����BŠI$�B�I�� VIJ1y� �q�e�C�I���X�U�d���ۥ`�1�\C�	�K[�| ��|��CH�,ߒC�Ɂ]�r)��
;�.u "(�mܺ�=�2gܕ+c�9*s�h�2I��h���S�? @�c7�_�*S��``M�_C$�ʵ"O�l��MSoJ�[��N�Z9^\�"O�����1���iR˼B�i"O���sk�:����԰x"O�
�,� /ӔбQ��1*e�T	�'��'ў��'�꽸%޵a,h�B� a���'4��	���1A#hSSAN7s(����'�愣�Z�����0k�$��'o��Ȅ��XQ
�C'&�>\�6�9�']2=��M��b������� ^~���'���7BE�b,4Hk�=q8P�b�'V�#A��VRMI�	�2p���<Y���������E*VUh0a]8x8��	X����TLr4�Q�A"Q��1rVE�%%D�L�@�Q,�6%��̃#,RL�Յ8D�l���9�N�a�^�=�"i�%5D��a/X�T6��;����\��o84��
�G�s�B�yFГ2�� `��l�<�0i�� ����/C��|�/	s�<!��
N�Lx��0]8|R�l��lΓ\�ڸ+���-��őB�#]��U����9a0���,�G e��ȓ����-��t���L�ȓo�©rW�Q��yYd(H�x�\A����?Q������]+�"J�Q�F@�g&�4�O��O"|b'�-I�j� ���O��lY�+H�<af&	�Mɖ��pN�B��B�N��T�IƤa2h��"�|��c���C4,��<$��2��B�Gb�R�C+�
5�ȓ:8M1n��[�*���X�L���$X��16
l����!���%�x��I&} )7�H�d�ޘK���dP�B�Ɇ:b�̺�d�L��b��ʓ�hOQ>�ӱƝ5#0��ǦJ�a�tœ%�$D����W=��1P%�H+b{���k?D�P��ܡlt��F��\��(�M(D��걍�:�ʨ�E)��`Z�h��1D���ƫ��4t�ʒD,�(	&*0D��!�+,hj���տ^QRa˅("4�pj�a5=�n����J O1��#Ѯ�d�<��.�3%老z3d�7S4�`7hMG�<�H�&<��!1U�X�Up�L�R�z�<���.URR	�&E�K�����k�<A�ɑ�LT��Pc��+.5����h�<�� �eY,����J6�~4�!/�dyb�)�':�~����$�4��	0j��ȓ'�8Yؼ��ً-V� � 	3�'`�hYW�	;7���
��`|��'�2��ţ^;��+\	ڂ��'�D�:'j��'���)��y�HHk�'��ؓK	8����(��01�'G�X�GT
%����М*��Y���	\~�
ˇwo��r�Z�P|$���c/�y�&�o�l]!ŗ#Bܝ�a-@��y⥑�"�h��ܝ|bmH�� >���0>�n��(��@Њ�x���,\b�<!aI�E��4K�T&����� X�<aU���ɂ��[7E;�����Z�<q����0"�-K3T��E����V�<i`����b�SpN��;>�D8c�G�<)A��/C�9�'T�n�.�B���ɟ�G{����.��p0���Т�R�a_j˓�0?IeDX<3Wm��"�x�����Iu�<	��NM�ç�y�v���AJr�<� =ِN<�J�c�_*B��=4"O�����4#kJ��1eԦeXV@r�|2�'^�ÈL
x���i�Q)�8�a�'�}��̞�/b\��@���	�$��'�ɫ��54��i��jO.������O5jdJT�.�������0N0���"O���"H�Y���6�ܱTAHA�"O|U�1�7�~�Aс�z��"OHX˕B���"���1s����"O���g��A�ɓ$��Pk"O~cWj�jg��j��ؓZy��*g�	Y��TJ@�w�V��Ӈ�z0 h+,�d>�S�'W9���b�')����V$�0�l����2v'�9�Ec6�^�,� T�ȓk-�� �`�;k�d�DeՈgK&(�ȓ:�JPAW�ټv�d�Q�蜇A���'�a~r��3�j<s�S�%�nQ��cX��hO~�O~b>�s�g	�?��A�&F�G��(#�&D�� ׇ^?p����7�Ϙq��YS�"D���Ɋ2s�pةGHM�$�����b!D�H+Vh̼W�^P�Cş?��p��<D����A���x����\�*�d���n:D�$�fa��m��,Q�EͣQ�4�ʶ�5D�$P�ц@o��IK��Vm�6�<Y�YK*l3��I5J+DaQ�(��<��>����B��q?��J!�?9��4��牡Y	ֹVcK4�$a(A�ȣ)C�I;`$Kb�G0:��$���`+
C�'�@T�b�1r��I=�C�I48 ��r�Ρ,PU�#탬%�ң=i�'H��<2���R ��cF��� b���|y��'�d�gĩ_�PS���F��
�ژ'�6P��FI/^Rz%K$,�������xb��\��9ӂ!�Cƌ%���	��y�O-9v�����C,�`B��y���
Jqqr��$TI��2KѸ�y��L�+���!�M���c�1�yR͋�I�K��l�X��!cP}�"��I��4�IK���"��Z ��94�¡H�~t���=D�l�&�G0J���a �B��q<�C�1�|L�C�[(/��1𓉃+,�`B�I;�P��`O8Z��M��H�/_NxC�IpʀAV�șH������޿S�nC��]q��١�$ʪ�dI(uʐB�ɉ���aoD��)0�	�d�xB�	�)� Lh��CƄ��1�*_aT�O��=�}����<m�by �J� T��j"JH�'*a���_��-�@k�Ep�b5Ŧ�yƀ��2H@+�1���A�=�y�O>~a��F��ր1�D�y�č�~, $H��^�$$�p�&i��y"�@��y �#��:��B�y��$UA��4��q�]r��@"�y¥ٿH���@�UɄ�Q���y�
јZ�f�k�	�|d�];��y2�X�]s�%��Y�x^��J��y���l�l�«H��Y���2�yRI�1""
\Zd���x]ܱ�a$�9���hOq��0{�d�(IʢQ�t�:>�1 "O����(``����� '����"ON���؇6(H�S,�6gg̉q�IG>�xeL\[�NW�#1����D6D��2�-L-7�h��b�_�Q�h 	#)D��p�b^�r��xӤ	_R��7l'D�� D\Y��]q@�B��5":ŋF"OV�P��J�u�Fa�f���U��`W"O�����Y+EF6i
� ��q9�"O�@��lZn�i�N�.M��"O��˦��],f$(V��,S��%��"On�ٖ��M2� ��K�D!;t"O���%��?��h���$Pj|`iV"O�iAbY�&b��	s������""Ox��vj�v��ÊF=gh�]h�"O�U��MTj(�̪+Y�Gd5r#]� E{��O���3 #�!�ȍ�UJ*j���_�g�ٲ��K�.�%O��y"#��hH�zW��<�V`1���.�y@�B�|�EH�9�r`� �3�y"��P���34�P�,p,���H���y��$o���s�Z{R�z�,��y��hri(�L��:��X���G��y҄P�s۠����5�bU�ʇ�y"�N�4���yV*�89V�x����y�hZ#Q�0p����+7�������yB�ۭo��xI�-�<��$�y�&��<ݑ#�+w�� �Â�y�!aR�6$շn�ᡴ���y�f\]�!����jXJ�9�����<��DѕY�����Bh�<�A%�w4!�d��(����e�H ��`!�d�Z��$�f��~ f�[�X�*w!��4�X!r��/�@�#4�	�!�D�?J<ޔ��	��<�!��!�DiL���l@VB1j���7Y�!��T�R�*�A��#:�����>v�!��Y�O�����P�fI,�f0Iw!�Ĝ7l'����A�&5�P�Ǭو{l!����zbو��ބ[N���eˆ�Ml!��o*&1���с?@M���~O!��+����&K R�y׉-.@�'E��i>E͓#n��#H݈N��) ��ץg�L��� V�i{��O�:����c�%*��d�'xB��6o�v�!�.�K�(H��Sc~�C��f|�X0��	Fӈ�Hp��B��qZ���`ǞI�>��C)6��C�~#�UA�F_�c&,R��N��C�	�&TtY��IӶ=�J|���A?6�B�	Nj���B��"D�nyQ�(ڗ99�̇��	u�V�3&�(�9�X{��e��eb&X�J��t��(Ϧ.p���ȓe���3�(q��������ȓeJr��V%V<�P�hV�C�̐��<�.e
��:s��(�АO��ɇ�]�	ƫ =�(3eS�G4$��/Q������#��9��̔��@}��Vjn��&"@!x��h�$��+j�X�ȓ%,���^(�:8Q��+vt*L��2J�kU�h�|a!�,�Ņ�]�5G^y;���G��FGؙ��Q��mP�� b-@�KG+��58�4�ȓ%VdB�nҪ;�0����Ev����irP�3"�Yڔ`�SO@%��4�ȓjp���ܡ��� ˧9+�H�ȓ}��r��9����a,_�O@�E�ȓ�l��d�Ap�SƆ��S�d��?��Dq��'yj�Xہ��n1��Lʴ8��1�0���؏\2�9�ȓF�͂2�:Ӳ0Sg,ޥB68-��S�? ���%	����1R���+�$ht"O "�L�!F���Ђ��m�h�"O�0B#���azs ʧp�!�"O�\���CM��P �)�X�"O�����7����Θ�B�ޜ�"O�h���_ i7©�̟'C���"Oj�k�b�($
.uw���O �6�|2�)�S?�vX����d<��hƥ*R>C�I3o�hX2����q{�Ɵ+"�NB��7�~��lS��]�Qa\"iTB�	��d�#�F�A�) XW-tC��KN��+�&��� N�B^hC�ɹ ΔB��K������i�p<C�ɗW?��jv�D
�X�Y��Ԗ~"�ʓ��?LOzu��+�}�3"ݭ:��Q��"Ob�AB��p�e �Hm���%"O�x�Dj͐`� @ba�Z���*O\
G�΅j%"J�$q|���',��ZB��;��۷�E�l��0�'Gh��w&�>Gu��A�hϧg�1��'=nm�@O�1�th���)^�:���'�"e�b�%y���	���8Uc��I�'q �#��$.�(�cr�K�l@�'p��I��
�h��T�&
<�P��'	3�<Du� H���Q��'$l��Ī,C�lKb�@�n>>�3�'Dm*e	L�I<����_�hp{�'� $c�
��
�^���U?���ъ�'ax�F�sl�
u-��c�f�;� ���y�L%��,P��_�p����yb���w�
mC��_�B�,�P'*�9�yNL@Q,�
v��j.(-ȵd��y�œ'7��m�h�.���hP��y�/%> p!P��\U*�*�g����xR�&lf��3%S�~�\�s����1]�IXy��'��MADY�&ތڕ���@�b�R�'�HjӇ�,}x���MQ1Wk����'�t�F�@�Y-
��䠆V>�I#�'P�	��Ĵ0��3%�Ήx!Fɒ	�'XJ���5��e�J�:d$Q	�'�&���O�r5XE���^�1�~4c�'�q��[/Y��.B|gZx�)O>����z��$'�M��dي�Y-7�'�ў�>A����ntHD��-טn^�9s�& D���d�=�>E8�� �qqN�� =D��c���=9��AR#��a�|��7�9D�P��@�z�Ȍ@��ؼT����53D���tm��1#4Q���-J��(*/D�|���1���)Ԅ�蝳�.4���C���!��퐤b#P�C!��\�	}���O�r]P1I��62d$a�퍨m�Dq���hO?�`��N�I�|qʣ�*NT�c�PT�<IT�	�����-X�Sc*�jfS�<�R�^�t��  ���Ōi�hf�<����R�E ����G�AB�N�v�<A��d`Ǖ	:P!P�t�<���s����	Z�v�>IA���p���Γ �2�9����Q�(�٥�9�Z��ȓd�H�Ag�Se�L��-K� ������4)���@:��4�
�x�6l��@z"<ICQWs���r��+e���ȓV8fx8��[3)޼�Qgȉ�Fj���CʸUC$O,#����>"h���B<�+�3a�4K�'��J�\A�U�S@�<� �HA�̌a|�d���[\��"O�]�$V
(�`J�jъe���i�"O9bC		S���C7K�tre�%"Oܝfc[>;�d=	��,'���%"O��[7i�&8�@u@�2j�J�3"O���ՉHK��)b��L��� ��D6�S�TIP'U`x4����<o�0Z�&O�'�b�|�ɽ0�F�A��Ǖ4$0���B�	�kϦ)i��^*U�e$J=(
��?�DB�-ɎDn�$
���Y��4P�.D���@Ҏ:���3�� �(��m-D�pJu�C^8$�k�g�16Z����-D�`���G9�H)�d�%*��l���+4�03p�ӌg�Ni-�B� ��f.�8�����`,Ǹ!�̩w@�j9֡�?a���䓶��e��J�C�Nj`�K�dנ0�� #D����L(L��)a��"�td��O D�8��
�$�hв@�X3Ṭ�4D�����h�5�p��$f@$	�N,D����L�H�����Zg1L�0��<��i<��c��/H�	G�A�M����	c~���*��q)@lܨ �ؑ� �8��(�O:K���
E�8�3�Z>Ld��I"O&�;#(�a�XPŠ�;(휙�'"Ox�ȕ�I�`B�J��K��ڳ"O�U�C@'�%C�D���ѩA"O�,�@��TB���Wi�:b"R�"O��+�`��.=�􇔴yTġ+B"O@�R��� i��tɑG�7b@�=r@"O���D��k�9`Ц�D�
�K��t>љ� ��uLx;c@�4�Nу� .D�����/R�~��I=?��x&!*D��Sc��C�����	#�8y�j;D�$RED�$E܄�C�6Z�0p%9ړ�0<��A�z�R,9�LH ��Y���s�<9�Ƴil��D�E�HD�q)�Js�<�#��+p�kw�S�6��tX���S��hO�'xd���%�7t$yI��,�ȓv��)p`�M���s��!*L~Ʉȓ���#�"�h�S�L��=0$݇ȓ�<iXp��!�<�PС��z�̇�n���G�Qw5^baOs�f�ȓ������<�aI�B��@�&���O��miTK�,�h!�-B�����@�'�f�s��r� Ȣ��+ZO����d,O�-[B-�x�*1��A��.�j��0"O��V�U`�v��`A��B�p��T"O�Y�Eѽ_?l=�&Mk���p�'+��a���Z科�95�ds&��U[�']a|�O:}|��pHN'��3ǧ��y���1A'��Q#�c����yRV vr�r�b�?�N�[�%Ԇ�y��*�X�ە�ȰHҘ�� �y�΃;���0�e�� c�[�.�2�yRg-!�YQȊ M��tA�[��y/�?���IwE32d"#.J��yn�:l�T�s��T?Z�� �Z��y"Kc#�r�a�9�%��]�yr��7GM�L�c�+T��pLZ(�hO���D�)�
�"��Pj�yrBP��!�d�$�8��]0d\�E��A�9^a!���a�R��E/$+�ȉf��<B!򤗮$���g��Nb "��\�A+!�$��D�D5X�@�Y�&�1.V*V�!�� �`�Ei��r7\ٺD��^5�	:��|2�)'m���@��>&U�H'���ȓDj�rqn�,{�l!3f*G�
ͅ�u�0MH@қY=$�(g��h�r��mv�ղ��^)�|�U�S+!����>cEk��U5O��̒!�U'T$���(e��k2M�`��"w��1������M=q¬����$쮅�ȓb�d<3	?�H� ��Q�v�j �'�a~R�}1x��猁+A�\5�ǋ��yr�#ͼ[beM�fH�����y2@��$�@
�R���q�K �����>� $x-lTL�L
;[�U�"OR$ё!F�H?"����q�Z4H5"O6�DkڶB\�[P�(.Kި�hO��B�h�j,ڣ�V����
bB5:!�$K&@��m����2\���0� �Z!��őgƅ���F{�VHP����U!�䜪3�n y�-ܱM�dq01�2C�!�_�"�ڇȏ�R�X{�cЏ%!�D8(�u����8����C�-c!�P5c�6�{3������?��$�dG{��$ERX�R���?��I����y�Q W�H���T?8��=ZEA�y�JE�i����b�ء-����d��y"	&H�@�9A�Y2�ܚ��L��y�F	i�f���\�vYL��'��+�y��ȕ{���	1M��? `�J�g��yBb�<N T eSgY�������y"#}�<���X�Y�vD�mզ�y��	Ln1�Ҧ̇Pv~=�q���y2�_�C$�vƜ=P�j�{",��y�MR�j8@`(�O��8�䋎�y��2G�r4��N�E�5Cf  �y��-+|V���I E�\���yBE4X���-۠=�<�ے�@��yR��!�Jy� ���;��r�㘸�hO���Ą��A9�C1$�ؐ�f�^�;�!��ʈ��٘��#:%`ݛ3U!�� ?	�)��.M�j��+8�!�D֫R~ ��$��O��Mqu�!�!�$�1
�l:��K����V�J�KR!򤛗ZǤ<cf�Y$��|�FhZ;)<��S���u����e�F%Yٕcx
CTD&D��Ӥ�C0O��(A
����	%D��H �Ɯ)k��1��(P���&=D�в� ��r�L �@� eLI���9D���J�8��M�q�6S��S�$D�8)v;]��#&N�Li��b'$D��QW��
KAj��Jit`SW�4D��{�͖
hF0��I&_J�Tx"�'D�t���4xD�(��*G'Y���Jt&D���wFͣY�v����h,����&D���ьEP��E:~�ąbe	!D�|�抃0v�`��3�M���>D�8��)4��\k�A^B���;D����%�*Q fu��#',^% �$$D����kH<i!v��
?B:����#D�p3�jL<}Ԧ�j�i�>n5"�:�H-D��t�c����� 9}Ւ�-,D�|;��8r]�� ��ґp���I)D��㏋�K��HpcN�<�T�.'D�Hc!��"T���(A���p�%�:D��� �oKj�y��]9g� *p�<D�� ���2�)2Z z«<"�h#"O$�Y ��?����� ��zU,�#�"Ol�Q�ǀ;��-"�/�_?�o<D��� �t�ꕩ	�TlB�Bs&6D�� C�I�ZCDH��*=b�(�(D����E��+�T���#����l$D��pWL.Rbn��E��o�R�yre6D�l�1���gz�)�D��|��*��2D�d����Dc�ɂ2�B�E��cц2D��s0���� ��RI��%D�D ���s֒�����5il �-8D��;�Gݑ��u�g\x�:|`08D� &�Դ=�tp�u��&Q�.��0�4D���WfAL�r5��K�<=-�C��m x�9���8ve��+�(*0�
C�	$C�Q�EM*��p�ң�33�B�I�
|�K���M�z�p��K�B�	B�ޜ���	mZ8S�f
X'C�	�];x3rȎ�>���B_�$��B�	n':�
 �Q9J�4�����B�I�8^@̹7�Мy� ��sD9v��B�qX���Wk_��[�+�A%�B�Ip�jS)�V��0����Hj�C�	  �����A�Q��6��C�I	X�8�fΫn�<hQw�]%1n�B�ɬ]7z܂��I�w�dJ!��7K�B�	)95
8�n	�B��=�r��T�lC��=����Ƈ 2L�=���[d$C䉻&�
!�	�Pn�Ud��Z�C�	"M���Y4%An�(�����$;l.B�I�Z]�9BW�=�$��m�#u,B�I�^dl�k���||D�BȪ9��C��I����5�id�.p�C�	�Y,�2�蔏H�>��6Ɔ�j#B�ɱvBȉ7o�`VbH;��Ax�B�ɴ HH
�.̝}�t!Af��X��B��[R� e�L�Ze��IxR|C��G4���/XV!	�f��nC�	.(�LMS��ޱ]>�a�D�x8�C�	�]���a9���Y�OA�Q� B�	� ���#߹z��9���&� B�I},4@C�،%4�	�����m��C䉧d�:�	��`��q��/�(c��C�I,T�x�p��a��*���)��C�IU���Qɟ�"��9��j� pv8C�ɕ��x`��(m��DY���+R�tC䉱k���p�ډ~o��qu		�B�,%�6�Q��W-¾4����jB�Ɉ&`L5��� �E�e�U�.&C�I/t&L(�UGF�"��M��Ɇ8,��B䉄H�X��բv��m�0��F/�B�	}vY��"�OD:ͲkF�  B䉰0D��WE�#7�JRC�Q�@N�B�ɥ;g}96/�<�P���O�h�,B�4t"����fd0�DF�7\B��3WQư�4��M�Ј��J�[��B�� ��ȓ'��uc�zE�&>�B�ɏ޴a�E%�E�F\�B�T��B�I�Rܖ��ůT1S�6�P	Q�6e�B��!y֤x��O\J"���'�tB�I�o\��20Z�)�ŐӉˮ84hB�I�c�����Z"�R��H6��C�ɹ��r� �q�Z�%0-��C�ɥJfx+S��q�h��NX�aѼC�)� �X�CF2o��l����}�F"O���-ފ�Fb݆)d��`"O�0k�A��Bi"�ǩV�(�R"OB��!��O�xoܐ{A��C"Ox����P�cb�K� 8w"O�8����-pf:uC'#�us���1"O쨙��e�n�2���9�����"Onͻ�a�X��%(����J�.��"OXh�h�,t�$(�F��VӌIb�"O촉�'
�2.�J�A�f(�a
"O�tj�%S*8 q@1�R'k�h�2"O�Dq���L�,ɳ�
OFj�|��"O�]�G���#��÷~^�-�"O��y�'M��Z��K1'��(T"O���������� ��h|*@q�"O����ԭv�>��h�:o]�r"O�4��6��8�T�%[��b�"O��R�㔋!L.���iØkM@)iA"O�	�F"֠t�9�'I2'��*�"O���f�
;��I��gњ!V�:�"O��2�`د!ì�AsdN=��Kq"O���IE�=�*A ���rx��"O�5�V'��iD��e"͵!�p})W"O8�
������0�� �?6�B��"O�HU��|�^���� 1��;w"Oɰ"^p��er0a$"� =�"O4�j��շa��A���OB����"O:wI�U���ZFM��d��KQ"O�����"���:4��h}tC#"O��L�*-���a�"AS��j "O$��1S5Q�.)��M����<ht"OĴbUł9DP0���>�VLS"O����u�F4a@Ȅ�	��y�"O%�W�$/,��9�	K�TY���`"Oh�⇆�)�D)�H�r5���q"O
1xS(�$��C �-BP�hs�"O�-8 D�?4�	�TG5��� w"O��"*OV�B���ۑ;a����"O�I��P<Wv\�eƞhI&x�"O*��A�V $yU�T�:���	�"O$ppv�9q5�h��K=(��z�"Oh����Q6���AIH�|��"O�uÔ���)�Q*���#�ru��"Ou�i}�|X#�l�=JjX�c"O$�(�qy8�[�{[ �q$"OhPY!�Z?,����T��;#�j���*OV)#3g�_���5�K5a�zh��'�f�J!1'0�$�U�Q\��"�'�8U�S��$)ϰлBkL�I(-)�'�J@Xw� ,�a0AG�
q�B�{�'wV�bEB
�OU4K0���;)����'�L�a ���i��2�����'�2,����:G��UR�(Ō5}��P�'�]��EZ�;=FaBU�]�.+�-��'}�m��J $e�,����),-��'z�(W'��D�� ���n��5H�'֦�3�F��F�ܕ3��O l����'��P(�'ē2�.�ꃇJ�c)�P�	�'K|xb�-�&z��q�h�W x0�	�'�d)xO��!�Zq�Z�3�(D��(P��")¡(]4k<9+�	#D���P�1'��p�V�~J�ւ D�4h�o�l��2�.�=�p� �/1D��p@�~� �VI��P�^�q�*D�� Je)�.��}LV�j#D\2FuZd"OJ��ܱ(�2�Y5CE�Z#�a��"O��!�Ȉ�{4Z�	�26#���"O����r�d��T��H��"O
q���S�}j��gڪ^���E"O��Ӳk�>U��� �u��h�"O6 I��,d4�e#A<3�J؃"O �H&��5�,8��_=Hx6U��"O�(��&�fVh�p�7>\
���"O(� ���,� �֎pJ��s"Oa	WI�j��%[ �O�%d>���"O�3D�[�|�֐
2GM61�̩�"Od��2W�~�)�Fƭ(z��!g"O`��K�=|Z�m�W��oW�0ʂ"O���0��*?b���G�N����"Ol����2h\x����lP�zb"O�Kc��,d����s��abC"O�a���u<N����6%HYa"O q���`B�Q_J.4�V��yB&̍u��%X������C��y�E��QS��g�X���R��y�Ƅ;%+�4:1ǣ]��y�/B��yB���L ��� cR�XR�)�y2f�[�PD��m^�in�����4�y2�_��Q%��mN0�!���y�A,
�Y��c���pGA2�y�X�h�.��r�N�=�M�-�y�jƫS�, ��<~Y*�	��V��y2���dѺ��!E0݈GE���y�nE%�\�[䇈U�܋��\��y҇�*�\d 0�ǧ��bu���yb,�Q������.DUt];U
��y�"��*�ꩋ��,C6�iT�Ƅ�yb�¤^j��H6�V-����DU�y""@�j����`��<	Z�C"Y��ye_!{h��J(1����h[��y��0_tXMI��2}�~U95���y����m�*��g�K�p����B���y"�U}~JU��;�<2D]2�y��ת��I���� 5��$�y2��VV6Qb�,�?
z0F$���y2fG=98�(R��P��qZ��'�yhM� d0� �Iڀ�+#���ybĐ (�Ĉ�L�5�8����.�y�B�	 ���3!,8�v@�'�y���?1����	Y6>���e$��y)׮Y�>`���`�,�A��yb��=\�
 I��1W��)jtGʍ�y��X�+xh���;R��C#Q��y"��5�(I�$`\t�uyv�ͧ�yB*L����2|�4�y ×��Py�M$��H��A�h,L£�]W�<�JP/7�pb�u;�u!��Q�<A�`��-nvUCDb��OC*DA�ONJ�<ѕi�5tmʉ�2lۄYF�I�JRH�<�iW�x���Y��8e���vd�Z�<�֫V�r&��3W��5Zת��E�{�<!���5PDI��6!Q� (��t�<Y�,<N˨}k��8x��H�K�<��̶�,��Á��θ��K�<�&A��>�-�����%�\��t:��t�Ӟ.zb �!JF�3.��ȓ7�%�L���	4o�"D����Q�R��b'��X$p��k�s�@��S�? ����珲���f+0�ڭ�"O@���K�Y��mr��4]���J�"O�ŀ�N�|��K"�:'�r!�"Oڕ��Ï�w`��5f}tL*�"O��{ŝf����3�U<^�pX�"O��-/�D@����M�z�8"ONI[AD�s.MX$�ܦp�"O�,�2��"`|{QB�!ȎJ0"O�ѻ���y�z�Z`�4�r�*�"O�d���^8�A�Q��gΚ�;'"O��kѤ�qC*�ل�_�PY�"Oh|��.�D5FŃ��	-�h��"O�8���]D�"l�f�@�j�"OJ�U*V�f"D W4t��+�"Oh���"X��DB͂e�F$��"O�Ei7@�}��U�C�m�
�"O*��4�רU<�q�@�jOz!�P"OZ�q�K[]>�t�p��*0��Ȅ"O�]�3�_'*O�� ��P�y�UB�"Op �O*�](�k =t�M��"O��0���.�,\���Vv8c"O�e�2N�f��]3�Mى(T�	J�"O�±m<�� �v���(Fz��'"O�	�t�T;hP�S�
B;KD�Q"�"O>��F}'�)���x$5��"OBIy�	J3�(��O�(-~��R"O�زNɸ`�,14(V�O^`h�"O���uO�%����'��7y�Y��"O�q�����Z��ď&kRX��"O�qqeFā'�m�b��"j�I3�"O
��#ᙩ*J.d)R^��E� "O�[3�Čq��R�M�)Ft�I "O�՛5K��:@����% ~B�KU"Otŉ���pn��%��>�F�"OjH�US�b����=z>Q��"O��� �?T�p��^�b�2#"O�(�D�Ԟ6�P8�`�^��	%"O����]�o���1�ܒy\�5�!"O`�d�1 "� �A�I��E#T"OF<���F���P@��!��X��"O��6.�91��`�7���\�Z�Z�"O�e����2oR�(!�`V�@=�3"O^��)_�3.�1)�6%[b	�`"Od)�5�α%�6@jFA�"v��l�"O�q�GB��u�j���V�ӧ"O�iT ]�"��&g��<��I��"Oj��'˘!-|
EA7憧5�0���"ObI���:Y� ��oU4T�ر2"OFQCFLƅ7z$�E�B�@�\�)�"O~a�� �Y�b��D�16�pq	E"O~���l����y��nB.9�ܡ��"O���B@�gatQ�l ���85"O�x1�ᒱ5m��0s�sl�ئ"O���f٫1l�JKt:Ċ"O거���
!(�%#CIϽB�҄!�"O����6@�"3��9o^`�9"O�4��J  ��p�pd� 1u�x�C"Oh�4�)1�=jW(X�'"O���f���&�4c�(Du�"O|���%Ȭ/����a�s�^$"O��Qf��z�D�$��6�K�"O��뒑 7�t:��	r��x��"O���R!vӲ�P���Q|tq�"OL<!�kŶ)\���MC�P�W"O� %2&�J�/]���f*��X��D�"O:- h@� f��b�� ���z�"O�0+� [��@�Z�hR�"Oց����N���4�U�LZ�ӱ"O$A��+`��<K���>M��@q"OJ�3�/D�>K���*C72��k�"O��cO�$J"a�c�$rZpБ"O�=ˀHݘb���Ð���+����"O�	�Qi�4ITk�j����s�"O�zR��:[�Pk���酨	!�� M��#W�NXB�))� !�$�g
\��кMB��3�/Hi!�_:a�" V��.//"��2E���!��RF4� �
�M&�5��	��!�D�:C�d	Ԇ�o$�W�'"�!�+e�	S��%{է��T!�һMK40�7䕢o��H���U$!�d�I��ű��"c��Жɒ�?D!�ă0|=෤P%N��tXdh�a4!�d��EA�yZ��)n�ޱ`�źE!�Ę�^, Q�m� �ɡ�FU>)!��T�HK
8a聳;��Q@�@�A!�D	�W4Nu*3��7/��hh�C�|_!�D&�4�3S�OI�h쫔"6�ў�ቜ
�p0�6�J��,C�v�C��&�������D^�R2ʌ�Cb��+��R��U�;��aK�b2�ڽIS�5�O\�z����A�(߶u�#�.g%z�ȓg�TT�%�$d�B�i�^�^���}GP���/P�%���A�Y:ꉄȓW�����  w��a�A"Q�1����=y����t�)+n��`Hڈt������y��\�XQ���lC0��͆�(O0��$�I.���4���9�p�BV	_���~]��z�	U���i��ՑR�
��1?D���$�X7��2��I93K�@S��;D��8H���WC�Dd��"�Y$2�!��
愴Z2�˲J��1�4\!�͗mxcU�BQ�tP�u�c�!�ׂ�*e�g�� ^�V�����!�Č�:��U��/��Il2aq��U�l�!�䋰|�^M��V�h���7�Ă	�!��%�6���O�M��(S�4R}�'��'E҈+��J���kHN8)'�$i���?�T��9A��ԃ��C80*6�����3��Io���%�SHѾ|x��k�2�2�/�O��PHr�x�b�.D��}��
���̅ȓ{/,���N
��9�!h�]�Jl�O<�=��X���J��V�V�v�B��@��2$���O���� �fm�<��'ؚ4'����c��A,�'f�'�ў֝�G���Cеs�P`��+vK(��D�>A@��O-��$s,С�FF�2�@"O:�#rπ��ժ�"��؆��l�OD��'/˼u���#ŀ2SӌŻ�O����0iYН��-Gw��<���ϯp=!�$K3y֥����®�?�j��E�����I A����R@T� ¶DacAQ-.�O6��$�ݦl��0="��A��G�p������)�B�I�@~pػg�C2l��i����!�<�>���h���5MB?�>�r�(ԀX��;�'+zUۀl��t��}�Sb[-�z�qT�2D���S���	�g.�.,M�=��/,O��<Ćs���Pd"Lu��j�A�<��CCD ���l�:����F�<� 6 {�+���v J�]�V�xc"O��rS<f�t�:3oA�!���Q�Oú�8U�0���zRa��>ny��'�$)YEjЕx�U8r�_��'�N=prȇ�\I��3b!P�Di��
���=9�a�q�V�5��I��oF��X�ȓT2\��C^�gm�l��Б?t��ȓ��j ��0Þc��[�I�d�ȓ�*��,>Ew\(��'M�>`��Dz�>!�r�²#|�TzF��6h��W�*��=)
�'X%���d'�M�L�1��'�,��H�ő�� �8'��6�D�'���ȓy�+��r�"���#r�����"O�Q��	�!IA���V勵�O���d�5��!А��.i�T������+$!����=�ao�)��c�ɑA�o~2��:��L<m�ZT�T��,��3� )4!��M�����SbҔ��1��f]t !���
i��\6r�����>M��D9�S�O�f�r�Gѽ3 v��2+	�$�K�'�
آI�}ڶX�q	�_��K�'gt#=E�$OQ�0��$�w���B�̹V�щ�'V���@%�"pP$KQN�^����H>����	�W�8��Ʉ�K5t���c�@2����w����O,��	�L�"��5+��8D���  C�֠	�Ge��b0�4���		7�	�'O�D���� ę�v�6C��	|��0��	-��h�lS$s�8B�5Y�T�S�J�l�p��W� B�I�!��t������cـ8��C�5iZQ�D�}E� ��#d�C�	�|r�D�' �&~��Xa�̱[WnC�I,ζ8��mF4q��%��>�B�ɱ~q�H�kU�;�pY*I-F�B�	=	��&*ݴtXT��bE�'�˓�0?1�IՈs,�X+7�ɍ�hdP���y�<��)7zzH�%C�p!z�p#Y��hO�O%L�xU���{I��Pp�Ɲ
�8�P
�'b:2@�/^���'�҆q�Tk�'����ԧu�ԸR��@��@�e�<��D�W�^� �͇�0]�T`�E� !�DS������7��Qj�`�!,h!�
���� 7&��.��Q�T�#e�{b�$ؠO�Bx1��F�D�)�Ĵ}!����4Ń��G�{.�<�r�,#`!�D�G%V�cjM�4L����-wc!�$��a�P��撙I}�e����wV!�ǀFҺ������.Y�����<+U!�D�����A*э?�:���*��H<!�d �����#�x��`ǌ�#!��OQ��@����aI�� >!�$�,2�hI��#J�0��H�4���ze!�D�.0���	�$F*>��(ժR�J�!�d�3^�&]ط���V~�tcƊ�49�!��0������tղ��7
!�$�2=4J%�F�\ t���':?!��V,����BƑ6#��x��d�
U!�$#-&�!�F��B�vY������O���Ĝ�A�d��ҨZ
|�)yQD�*|T!�DҚ[v�d�bn�Ho����b^���'�ў�|jZ�=G���4���*�A���t�<I��)x7�}�%�A�"┑���4����tI��6�p`q��q6���IkqO��P��%5����K!u�p$�"O� l����"y�΁V �'�JR��_�\���A	L@ZaQHB��q��#D�t��&O�&0y��۳�$����"�;���D�1� �b�D 'a���3Zh����<H�,�R�.˽#�dҷ�#D�P�eˮ��x`��&,Mp��N"����Y�O~�P:t�@�Z�̖�c�w�<�ᤚ�I� l��h�OqB�r�M�r}Rb�F �'��i*�Hi�yQf�ւY� ��3k�'hx#?9'�ф``f�F�An�RE���9}��۶�i��D*�OX<�I�F��Įǣo�<����'��O8��|�M|��
������%� j�	3��j��B�ɩ���-D�.&���RO�.|7-8�	x?�~�,O��B�T���&��O�2�q"O(��P��� ��6��7.9xa�B�IuX��P ��1K��\�Qꐲ;�C�f.D��Q��#�u#qE|	CP�ΩY!�$�^Lh�SJpX�%��U�!�ď/yV�xdƈ:�(�Pc
�6)�!��A�b�\��&g���C�(ф(�!�D�+da��Sv�Є.~H<{gW�9'�R4O&�0��R*�
��VG�!���3B�����	B	��_�.r���D�H�">�S+'���m��[�%��y��L����y�A�+it,K�g�jCPP�����OP#~z�H@�@'�Uib�2Np֜"�DZ�<ɗ#��Q���aBQ�e�(�굅Y�<q7��?Q��d���%Z����Q�<	g ��_��h��K�n0������P�<if(�"@ �Sg�A�]Ʉ�ѥ�I�<�DE�%a@��z�/I� �:��GA�E�<y�jH�h2�XR&��{b���#��}�<����rm4�:��#}1��0�,r�<�p��[+�2�KР[�Ѣ�Jf�<���B]׬���o
�V�d����Aw�<A��״*���BL�r"����Po�<16'�(��4�0H΅����Glo�<�#i��Y>е�/Q�*�fQ��RE�<A0�G��d1W�ۛY����!��f�<���E|�ܢ�O�>w�J��b�<y��Y�@EHu�#�:3�ཡ� PW�<q�D�Iu>�+4e.*�h�ѳFUV�<��!M���(�2H(a���Q�<�b�t�.���H�E������RJ�<�&@ߡY�NXXTCR�cy(""nB`�<yë�^��T9��'IN�u��GDV�<���0�z]�f��p]nQ�CV�<����n96M�C�L��(^F�<�B�Ctm\��,!SXXDx`KE�<���F(`0��0jM��z�<	2���4�rdș,+F��A^y�<�0�#[Z���E��G�FDP�v�<��P�t����'�,_��iy�(�I�<�ց=E�"��s�*z�`A���C�<��`�Rp<!Q!�$�Q�-WW�<Y6��Ɯ��+��^����n�\�<q��8�͋�'=���B��\�<I�E�-| 0���;:�&�Y�lD�<1p���^ =��b�5,��A{���vh\\:RY��K��X|��Z�KK�4p�)D����,ڂ�G�Y�A�ƴÑb$D��q�-���"��@i�%������$D����ȓ� 0@���OПZ�BEе�'D��l��TXi:ԦϜI2B��8D�� � S	0e��t!�Ȥ7r�I�"O��錆o�|�i �í}����D"O��B�,}}rU�!��9��q��"OL���<N�N8��T9�H��"O�hc�2z��i�ug��N��)�"O"4�K(L�l���h΋��H�"O�x�"�A-��A�fY���ԡ"O �����L�➹v�	��"Omy��,uL��#�!�3N�,i�"O�ՠ1cμo�JP ��ψ ��DI�"O����]>m$�� ���US�@K�"OT8UH���h ���0uA�$S"O�-*��G�<<{�M�'5Զ頱"O6�Z�΄�_�\1Q��ckJl� "O�q+į�CP0���Ss l(""OJ8�7�$�T���/�:o6	��"O<T�#�!</���"L�V=���"O�ѥ��v0̳a��Q��4Q�"O��R@�/n��d"�kD�i.��kS"O<=SE�U0r@=����1�����"O.y0@G�#}2����4h�<t0�"O$�:&
h� 8�&e��n�x�!"O���ȟj��5��dG�
$�z�"O𼢲`Vz�H;��=�qb�"O4EI�B�"	�@(��d��M��c�"O��	P���O���Qv�T�1"O�YId�ق*~�94!ի1��P�"O0�Շh���1a�D�<�Y�"OjI ��N�b��	�`�	y�6��"O��z ���8�$��p��p S"O��jq�\#����F\Ox�EX�"O��⋾��x
�R�'�tP�"O�x��iA�b�c��M� @Y�"O�9{WfJ�v*<��ELP$��99�"O>\�WޙM�	iA*�s��;�"O��ɱ�_02�v�s��׀D`�3�"Of5���]�N��V�[�/�v��`"O��#��1P�tH��Q�b�X�`%"OJ\����j>IQ�!F�;�x�i�"O>L�ѮC�>R8�BSd�u��"O`�h�$�!X(x�P�A��,V&)×"OY2Pm�p;���� ,N Y�"O8����߲tG�<�<s)@�  "O�i�o��My⌑@E�B���'"O.]b����z5)2�Sc*����"O�%��ۼZ��@e	W�G=�5�"O:�`�Yg ��t/�T,r+v"O��	6lH�|�A�)۰[~lSA�'>������a����!�H%-Rt�;$��IP��R�'bj�I�]*+�l�3��9(n�-ێ�D�Xw�TJ��*§Y��s���L�)��
ψl$����	l@-��'�7r�<�C��B��poZ�����6�߆C��S��M�t��&�(��T��&+�Rm�t+�{�<���IJ���K�y��D*��v}rnV�[�ħ�Ix�8��&A7�|�ѭH��}D`6�O�¦�/a��08Q�B�Sp��t%
en(����B���x"���!�E�岑#sK��HOj��!�FÊ�4����UP�B��U�`[)�y��S�Qوd!S��u��10e��M{dʛ�*hr`�.?}���iʌ���g���`gfT�V�����'ֆ� E���k�ѺgI/G`QЪOpLw�W?N�t)�d��C��g~��0d��Ϡ���!!"�]�K��Rr'+u%�,�(	�KL���'q�����b���g@�3lN�Ӎ�dל�Ů��>� x$X� ;.sh�k��9am�T@3��d
ĸ�"�'����MJH���Ç""8�\��'ޠ��ɝ��|��n_��A-O,�
ь�(���7  �v���"O(!pԯ���%�HT�� 4�|2N�KS��0d�RB�O	��i�R��}ZF��L���pD�9p�R��%��U��9)�D���~�B �J���	=#��x�O��w%�	>0�'��ĘP��!r��m 0`Q�6�!��'SfX��$<O��l[�X�V����.YNv�D�*ɺy���E.a��!V�c?m���#s��h�&���d� 5�2O��c#��$�U:�L�>Ѳ���p�|X�N�'!&�z0��;/	�NF@8YT M���g�Kͮ���&X�t"��Dz�\�O���@���6�<ip擑]���$eݚ�z�A,5��]P��4��X:�!_�!+�B�Fq
i{@!"h��]���]�9h*�3����	�g��	�I]�æ`�B� Ƀ��:+y�hB�w����&�2�� `e,T�/
(���'�LQ���4vC�!K�`_8b10����2�(h#W��3G�C�C�L���n��#��"��4�Sj}��ĀJST8���rA�����p<A�d�_6�u D�H}rɋ
bx����h����^����`��#fX��N�YWJ��J[�'� ���F]�r�h�ѡ�ƕm��O�Ԃ��(4�<��_���4�[8��@� �>T��d���P�V�輩r-�8�,�@�=:<A{%�'��X7-SO���r��ӫ
���q �	��Hm�`M�4W��Nڦ6�\�Ū�'W.hR=ﴝyâ	U�� K��ݾi`n�RqOZ\j��!FjeM䦰��nB�a6�z��1� i!`J�k�>Tzƃ����ST~B�E<N	�U�#��2�t�(�&��x��T�"�6
�oUA�-R�a��D�i")Ң$�)���2\�L�"��1$��z�� ����&��B�F���ę�Q3��1�k܅R������F�!򄕌{�
KT�O�B�\����/�1O^�9V#Ə-�Z���G��!j���t$4@@o��+I<`$�72�a2eA8r`�|��A$D�x�=рB2�gyRLF+�H�ƌ��r�ej���'� "=����B4�L�`)l�9�3%1��3"O2�J�^�Qq�f�D�	+��0"O~h9 Ȍ=i���e!�>6��"O@=��!INi�QڢAH�I��0"O�13�"|Lm�DO��Q"��'7�'�a�#LƤcp�����()	�'>�-��2:D��Ə��k�A��$2?�S�]�n���p@��&G8x��j,ݬ7~�i�"O2-�U�#�n����Wo�8P{T�>�/݈}�ֈ*�-�Qė~~]aFlҐ0_���"O��ke�	.(�fT�#���C7� ��9W$����Q����	��g�Y�8ɳ��"G҄;�ԍ*d����ɓ��a�������-JXS�R�\�����9}��ń�	�g\����/6����T�5*�p����Hk'��51ktYqU�^�
>h���~����^�T�BuX�e��XY8E"OƑP�ٛ^�`q�捐G6���O��'�*5g��0�^�o�N �\w��Ɋ�����o�|�9�&���PK���p?Y��ϟܱ$�W(V���[�q���%��Oe��P�"�k���)�m]�U�~���'�x��)�]���P��j��pS��D�%O@�'��|{�m�O ��]6�By��aB�5dX١ ~+�EkA�T7)�{�kѩ*���s)ʡ��q k�6݈O~!�וy$4uY��3h����� �Ǣu�vMrC�U-L"(��E~�<���@ht%��-^d
ђ�B�<���Y��� �aQ.o&@a�A �8@i�Vw�a�@�E
�_tfMX��W��q��I�W���	 9�X���,
�:f�I�.1�1��D�Τ`�#�_�EE~���C9�d��"�TK`)�b�<���A��0�a~2.P�X�=����]���ːaO�B��`s"�������1	��1lO�8q�B�D���h�e�#%^`�R�>���>14c�$� �jf#\f��H�!�%C1JT"�H���\�R�$ɍ<�B���lH%3���!�'j��
b_�iiF[!#�|i��	!#���F�38�d�5�F6��?^�ؘ ���T��D��U��"E1�0��r$�!�y���6�a�ËFt@t ��qRNl��H �4�pd'D�%!dAO?}`�(�	LN�2�>O��ɢ+�蝀�ꜦW9�t��'��	7(�
�vlނi�Tܡ�\6u�Lq2�|����Oi��iCJ�&'�,�l߀m��� ĕ��e�� �JB)�`�v��e��<��倐��r2�.b�~��E�*S��)$D�=H^�YM��wH���j�DNp����'���!)�9���v��1,�*�B�Oѝ�ā� jB�	�b�U���q�@?����D�0-�.�R�Oq��9TFC3f��'A^�"/ޥ8�B0D��9q��
eB ����y�E��T$P`NP&Nl(!n_��!�B�� qjP����i����5��V�B�(�u`E��|�����d1�Ӻ3��Kgo��ʦK���J�˕-���b�� R�rA����$a�R��A���-�X  �
�&l�eR��U����S���Ҕ]�Y'�V'$B������u�+`H3}���ʛ`�� G���S"+���`�}���&#��B&��B�2�
h��lSӣ�!g��a�z�2��CG��mڡ�Ox��U�b�)!�W�k�R%;�Ў*"e{%k�Nli�V�OtPm��|"i�X1'jP/:]%��, R�AǏ�D�.I���4����48��D{�;k�j6�P+4�=��$�eY��!dd�:s��N���q�Pg�,6&�(3�%�������>'Q ���Kz��9��Ō��=���TD���b��$���ȷ4�:}[� U8`&���BO���L+��6gR�v"�O�����'��%J#�˙O��d��	=^�(�O<��'��Iҗ��@olqE��(M��,���/I�>p�i�F@R�K���	��$����l  ��¥Ҡ��!�P)�TIb/n3$HzQ�.W���y"S?͐r�Om�(�e׶$��F*��i�[h�(��	6JS��:	�'�,E!3���l������Kl�Ј�/[6H�"9��l����fH*��a�odPA{!ԥ�?�/O��$@B ������5C�D4st�#<�F�K��rE�k�4{��I�k�� ����$R���?������%�Nȣ��ik������'
�"}R�&ŁU+Bea"��'��� �TjX`��u&�r��`� %făV/Fai�/��	u����x�Hx�O�1ɠ鲠H5D�P��BM3:��'�yN�Ke�G4K%�!�|�n��'��Oz�	M;.�я}C��L2��uK�:[�j��`GĴ��=�J�	z\|렣��M�pT��+�M�4ض�>l���)�L�����n\���x��xC����h#�ʞ���?AЁB5~���&��*�?��?>T�W/Po�&�2(� ��5s)M�B0HM��'AtIx$H�Y��Y#B�<��h�B��A�,����4�?��-�$,K`iHd#�Լ��"�/;�B���ʛ�vxc��	W�<��a/�`b!�ϩX!c���:Ij����#Y�������-�p)2��F+P�Y[&���LiB���vp��'8"��ٮX�ݱ�jT��t 㢇K�.�x��Ѣ
$*8-Γ.x� �rǻ��=9b�TL��AG&�H�M��B]�e���G�8)wX9�O�%�������k[>~�ެ{�*�o���*t�y2-�7x������*ZIj��P���p�w!_;_��O�|�G�s�ų�'�L�2��7+�CCd����;�����SAJhq�%W�1�� Lm���`�*�<�ӫԚxO<�$G�~�:T����}��qЂ��Mh<��W?D��*YY�4)㡊ğ�M��H�U�`%#�O����W2{m���AL��W�*#�}az��N�!x�����bHˆ���^[���O�����R�KJ�y�f���x�=	�%�����cGȐW�]��8SQLE�MŲ���@��I}����"sѢ�Ȳq�����I�
��'Oĩ�%)�[��yq�`��h�1���oN�7M�q���+㊛	[��UPV*�_�� Q���r�Ot�Rc 8�����J`PX8�'%��g	N�%�P�a��K�@�s�'@v��S�	2K=�TN��<A
�'��<�v�ԯ	N��A�eZ���
�"O�C4�ا_Cꐱч�:���""ORM���	Or=a��Y��W8�y2.�@�|	(�FN�M �h�J�y��ɇT"�B��C���q��)�y�
ݹjxH�q!F�GzQ��d�y��&:�����$�-;���E`�;�y҄�w!P���p=��#��y�霃gT����_�e��,���y�O�L���.K��X�t���y���bL�����ۂ��c`��y�o�. m�S�O�yC�<a��M�y߽]�@�q�.�3rH�4Ȃɖ-�yB�H!F}h!�\�w'���CT�y
� ���G!�T�1��(���8"Ol]���ݙ!�|9�C�]�@"O��C���c;����¦ j@Kr"Od��Ճ�2q��

FT�"O���3$ܭJ����jȳq؆��%"O�
��ԷA	� P�IZ����f"OD4B�퓔m�@0�^���%c"O�ak1&�A�U���]N��JS"O��#�	C#����dE4)��
$"O�]cf��(��q��B��V�<İ�"OX��R���0�<
��Tz��%(f"Oh��F��pC�BߨP����"O�0[�AL/p��1"2(Y��b"O�bQ������A�W�P�Ă�"O�`�A�Z�G4�5��`?�xx"O���Aַ8��� 7�V����C�"O����H!Xt�����_⪽y�"O����䞉==
�)֜�\�Ц"O���CĔ��&b�4ղ	%"O��7�7sl�r���=S��s�"O8�ۥN[�N|�� L�`@<�y�"O������M�y��Q-6~\��"O II3=D�ha�hѲ��e�e"O.�� ȫ)�t�1�Ϟ0p���"OL�d
N��"�+XL�q"O܋TԳ ���+�E*p��I�"O���oA;!�t�A�ARؐ�V"O @� �H�[��0��ɻQ��u"O��C�Fǯe�z�Q�C>�P�p2"O"a�V��1]���
���+p�����"O��BrF�T���P�	½ �!"O�(�ԂFF�2�(�U��a�"OH8ɶ或��@	���8S�09�"O���ri�[<&�{��̵��u�'"O�L2A� � ���2%{�Di�B"O�h��@�zxP�a�)[J�,��"O�X�v� �88]j�S?:<��"O ���ԉi����ӑ/҅�G"O�	q�D	"�x��'Ѿi ��Ҵ"O�tI��O<F��̀c���x��J"OAb$ǝ��̐�f ���;�"OlpZ�A�1AML�q��_3��"OF��`�{�D0�ф,F};�"Of$:��&;+���!� �t�h�c�"O�%Y�F�=8稠�w#Z��M��"O�h� �еU5�lC4Oٱs��1�"O�����YQ"���wo�)��ݡ3"O�]`���#'���*͞���h�`"O�t��"_!*ĸ���2�f��R"O�}bS5VJR�Q$K��d�3"Oj�PM�OH�ȁ��H+��Q"O$h���x]P|r�n� ���'NQ�� ~��|�Q�/N�4��s�ś2Y`h��'�dձ��ω}���#C�0"�"չ��Ď.[pf��SB?§5��"�hH�Rx��⛌z���ȓ	$.���@�	֤UѢ�6!{Ѐl�W3��Cڵ+[�S��M����]�$�4�?/�-CV+JQ�<a�˕&��LY,�7�dX��dGS}��Jd���8DCex��@��`x�P+d�ܡFh ds� �O��F����{FeV�t�*}�����KrQ�jʂ��x�a�<.Q�Q*T�L("ȋ�AX��HO����ߔ.�&���$�&)�
��9/��;b ��y�-����S�ٻT�>�0�ʒ��M����0s2C�j0}���i���с+/K|@Jࣟ$<��\"��� �){t�'	��}����"H���1W�@ f�RbfYʄ�'�̅hr��y n��u�H�]��
�4�*1�8O�=�2⌕��x
Uk�f�� ���:4����&�1]6f}y�镹?�9ƫ.�:#�a �����鍡P���@�N�$I�B`���;a��5�'Ud���J���(���c
�l�,ț'����PȂN��|2dᇮV�l�(ORy�IƱR7���r�ӣc�0=�T"O�H�ÎN=�XJ�qD��H'�|
� rC��xw��d�O���#d'������r�h�h�GPCt�����:��Ĳ�K�	R���PH�	���	�-i��ɸ4c�O�~YjؼV�'��y���>��YD���
�j�'��(a�ʝ"/��Y
"�;HJx��L� e����$&����dĆ_��H$Fb?U8�%&@���M�Z蕠��.Ox�01&O5_PpM�¾>��)e�.d�g�Fs�FM���Э+3���ʠ�֣��gܓ0k
�KG��G�T8X�%Ą_RͦO��H�J��� �E&�<i��A�-#$�)6��q����D�S�!��y5x��E�A0D����I(i�`슣u�dq���ɡz �ԁ�����'O
ᘳH��Ä!XA��ڦ��@=�<B�w�>�x�C7c��BwJ�r暱j�'p �&'�$YN���L�o�̨a��.mym�E!T������@1F��槐'\B�Зܟdܘ�O�p$�Ge�!{��
4#�İ��'���&�H�/^؄�O`�1�j�4*^`	�Ȓ�Apb��Q,�q���#"�q�(�+�g�.����W��P��WD�L�8���Ș%�6�iXW��3Iʓ#��LE�,q��n�D����$�"�[�|afH�7��:����dV�YK�D���\�O�	�栍� �n���O��+���N���Ywx&���D�&�Lc�f�y�M\NQ:�ώRjݹt>��x�kǒb2E�Ra{85!���|jivÑ��� ���*�hr$9ct�i%?1���k�D%�7aa3����f^��xC�P�PdB4���}n0H��͠g�@eO�$@�pa��	�x�L����d��0a�Q�����X�f��m�����Q�)�p�`^�@[.�s�@�_!�ĚQLX%�b�.0�2D�E�"�1O�H� ����E��,6@B6@
H�Y���g�<��+؛.z�C�h�U<(�������=��.�gy�J�f�>Ab����y1����ʜ1�y2"uA��`ʛr8��{��)�y��#�Eũ	�aV0�0QCQ	�yr�Z�J��Y�6���\d�ؠ�ߙ�'8P�� fT�/��q%�Z�p֮`		�'���x�+�1|h@�m��c�����'aY�K�t����b��T�P�'N �[��\��m�S瑟l�
�' ��pJϋp��k�&�,l��
�'��p)�*G]<lRajU5x��i
�'v�caO��FMX��`�K ʚK�<	��گ5���HH�f�����D�<�!(ã0e2�i�M\8E�����@�n�<�ŨA6Sul���4-�̍s�O�d�<q���^Z �)T��0PO|�С�Wb�<�C��c�� �7�kHY�<A��O˺|u/��S��UP6E[�<qs��Q,�8ЬS2,�j�b�l�R�<��=���;&�,�T$Yd L�<�3���Y��s�(]-7��(�+J�<Q��E&$���A�\ !RЕ0`F@|�<1GĄ&�V9v�ȟZ�
9�&��U�<q�E�T,1#2�գ3�rI��M�<IwN�=�P,���L5��Aco�S�<��*�,q6�*��Z�B�󷋐g�<	t��3Ut]�qH�2���j�o�]�<����i'���M�Z�rͰ%T�<�P��8>�Nt�G"��,�٦R�<���;3��(@J�)z�ցYR.�R(<�u�]�X�,`�a,K�C�R�6G^�o�N̘�����?	@�X!�<����	z��̇N��AF��\N\��>� �"�` )N\�(g�D��U�"O���0��F�(�R�&,�aA�_������<���;�E>�sw��=$�P��@�|l�B�;D�XeM�#��Dh��"*0�S��RҀ˓TN��� ϯ��g�e��1��JI}	LR����e��Ɇg���P�E�8�Qs���p�M[0%��F$�3A�u��@�VgɄk���� � A����kw�D�6�!�i�%� m�4�KT�[�#=�Гb��6�x�Ɖ�RP��`MJ57���"O,ر$�ɲ-������8mɀ|R�<O�$���8Y3佳VL	�'�$̙t@�2/�����?�ɘ�S�|��)Xh-�(���H*&��{�ͣ邸R�����aʧ�ԋ�����.�⽚���@�`� ]J��زl_�L�D���c����A�-�8�|����Ѱ&E�O,*V�	>x(Ȓ��D޿PX�4
�Q�t���M�~�88G�E�I�M1�K�
Ԕ9�W�'���S���F���bV��l�ޅPV([9C���Y�I)}�<��]��hS�U�BY�Mи�eS�hތmq�<I ^�< x�2���;�!�d��	2`�̿6�u[�j��� ]!Z��+��Z��r1��*���	J�Eͼ3�}'>��ݷ`��8��e`9���0|O�59v��09��
۴kp>E�ā���t��7!�{L�&G��J0����G}���OR�S� �-`�d| r��\��5����R�e�d��'���H�P8��
�
&�9z$�\=.�V�O�E ��P!d��`	��49hCط.b�K�$�%�Rز�S5c�i�2�>����dR�&�\���Ӄt��PI����)U�G�V���	-8�J�k�T�	�#v�-z��ƛu��S�D�$("g�#Umh��&��������S���NK�X8�X>
*urg ��OL����*�8���'8@ڔ.��:rݭ;+�@)G�F�f�a85��doRH�I�sfn|{f���V����L����ȓ�%���{Eл|�B�������z�HʿS��Ӈ��~�=)D$E#(5����E��l�Ve?D� YT���|�	Z�FH�@g�ZFO�ؚW�[�qg����J�O��鎮�!
�}�BP�Vz��B��$/9�Ð#���=��#>
5ZY���Wt�$2�L�=;M����rk:�����@�CcQ&lI����ԒVm�A��B�O(����.�:��O�hgaS�#��P��O�OT�3��\s �JZw�D��DX���+�a]�h�'2fy���22eJ��F��5%�u��\,�C�F�<�?I��+\8rY�E�<��㗉΋aQY��	ЁFb� ��,F�<9�F߉/�PT(#d�8t��!ʍ�Rn���B˄�6I��C!�џ��S�-�@|x��$�5&����¹F׮�A6	��{b��g$~�����4'����	�b�E��,C$��c<Ob�q&�Ì���]�a�N�$+(	��d���]��� ��: Ǝ��X��D��\��i�0g�Q���)p���c�t�!���*)�XL[���rV5�baW��n����E��,�%�"~�ɥq���n�1'��8����adzC��I5"m��MI;"��P�/� cTTC�I�;Pu�qJ��hm����dѨPFB�5eWA!ڱw֔�&h�j�NB��(�v��c�<"������.B�I8/
I ��Q"F�ъrh� !2B�	�ں��]X�J��oY���2'2D���q	ǠL�Y�ꋨa�	j��?D���c���a\� Dh�EN<D�*4
P,d�}��VhpR�;D���Ԋ����D q���r�9D�D0E"ɱ5����#6�1� 5D�|;��ȵ j�:�� �3Έ9�O5D�ܘ���XԖ�Z��#:D��AJ,D���`�Z:G��%(Į�R�p��%o9D�(�2��@\���ÁP�tT��9D������*'T�9��	���!eb6D����)(A�� 2k�g���2�7D��J5��<<y2Æ�J�Խ�j3D�P@�.�%�\��!λ,솱���1D��
@"R4m��xr�A�G�|I��m)D��X��ծD-l9x7��#U�K� D���C�H�
�&��B�Z�jZ,���>D���
�!�,�" �M@ ���:D�� l:T$d�"��/LH8X �q"O�40�hɝ�5���Bs!�I��"OJ-���T9}���IQ��8P �'������x.��aK��Ob���*�"�S
�'�Vl�wJuɔar0��;0�B��	�'�<��W��p�βRA��R
�'�@d��Ǌ�V��99 ��S�B�#�'uv�xb&=C�� " \�G�� �'�^�0�ޏQn�B#ښ=�4���'E~�#�ٻo������D�)�'��l0���:�%HS�Ar�@��'�Z 1�F�@��鲳�G(&@5 �'��!1�Z�Zy �\��6$��'���R���fg� ���/Np��'�R��D5
i8mp��I�3`hj�'F���)ّA�(1k6�@�   �'.`<�tm&��ي`�"^�P#�"&�S��?9�韚
�,�%n�y}��Z0�j�d��z����{��4��-08~t�S�Ϊiφ�Ѓ$@�~�CrvTI�=�O΄OntKև��%�Լ�RlI�c�����7d|�SBn��(Ĕ�S�Ĵ���?�YG!�Zȼ�0��U��lA��u�t���ۏ3[X����`���)ݢLV�Іd
�
����	���)�4a��mI��`��!K����O�bȫ�I_�"���y���d>��)O��3��&gV��T'����n����(�7�\A@�#�	 t�r�cADI�)�'X��Apc	�/_��ɓ"�K�g�d�I�7����E��|�)�'E#��ca��>���s���9��TY$�ظw�5���@�
�'L�"��?��LS�,�r�:�:Ф�-l�<��'�����Iu>�`�� c�~ݨt�G��H�D�G�8��8��w�l�Hp�V�I����?٠�4���M����9|r�ȫ
��9���CC�<1� �!r��+r�"�Wo�D�<���h���j�cX.c�x-k7i�B�<A��Z��3�g�4=�0�*S�
V�<န�_�j�!q쏴eT���0��O�<�w�:OH�zU��r�ԑ�BK�U�<�!�U��@Ł�Di��@:W)�V�<I��5;(���!�N�a���ѳ�]~�<�BFߌ$Q1f��{5~|�OT�<�� {���8�X)OqDDN�<)���an.�2hO�1.*1q��E�<Au.փ+zEpC#��qX>!��E~�<)��A0V�Fa(�gY!�r��a�u�<Qv)��<`�b��.�nب�d�s�<�'��'Z.����)�:Q+# s�<��G�_.n�9㩄�|јŸ��G�<�'-ht��S�[e�R�p��G�<�Uᙬ47�5-~�x�DX�S?l ��H4�Ǒ�R���0ȕl584����hhP���1� �FNS�:K谆�_^�����w)����m&씆ȓ:�ؐJͅ�`V�g@�=�V	��:�P�`������h�cfՅ[R: ��{&��7��GOt6F^�f��M�ȓ2�0ӄg�Oà �S3�~x�ȓoP�5��@� �ba!�zm ���r, �Vt�A��F[=h��)�ȓذሃm������%�>E��mu�i�䮇�M^Й�k��#�la�ȓ\KTй ,�9j�� $�:R+�<�ȓ�&A`t�Op[r9����0<��ȓI\���̄����H���)L�I��4��8:si�&�]��"��@F�Y�ȓ.|�h�EjBc̽s�N�"U:!�ȓ}��`��k
@Jx�ԞRȂ��ȓQP�	��H��=C����#d@��S�? ���%$2Y���#ċʬw`쥹G"O�|S'�U?����Ɖ?=隕�"O%@0��Z���b�ȉ�l�)b7"Ov��E��A�0��hǳrj���C"O�a{�����0"�PxQ>��"O^u��o�"��9�$�YC�i�""OT��@_.Rl� ���h����"O��%�ji�s%L��d�z�$"O��@G̘�xH\���m�6C����"O��s`�ިTp$���̀ 7XLlä"O�u[�G=^��$�:O�f��0"O��[d��d�z3���R/�}`�"Oı��E��8
��铯Q�r,`�P�"OĨ���<q���-[8�pܚA"OHa�C�5(_nQ�D.ǆp�T"O6i9e�ŨB5��K�N�k�"OВŬW���4R��R��U�3"OJ9Q�� ߨX�Ɓ�}�p�(`"O�ZP�
pXn��&���>�R"O�L�bk�y��2WĎ�y��yd"O�� Qg����X'mZ5p��\�"Ob��!W�A���\�B��"O�h����/Aw�ctaQ�o��ҁ"O�D��a^���"`Yk�RS�"O���R�[� O�!D���"OD�A�͍@��� 5�V	k�6X3"Oށ�$�7!��)i���K��r�"OlL�V���=� c�5u�ɐ�"O�t@���(爹��g�G���!"O�I;eI�N^�}�6	O?35^��"Ov)��H�!V���@u(�6*b���y��֖>�p��ȈJ	�@y����y�D��m%V�pA)�:���s���'�y��l���૞ �<!�I�yB�X�5GK�hwQȰ���|هȓ����S@��xX�! �� "-���$��#r_18/��c!�����"D�L�W�\���鐩Z4���5�!D�P�ᢟ�m�@���	�)vH4D�`i�4T��Y�G [�4� ��'�2D�P���"vah��Qn�Z0̪dB2D��ZpLE&	o��@ƃ���<����1D�+6-V�slY�4xjtb��:D���i:g�� �k;Q���6D��
p�D�}ꀅÔi��+Z�2�)D�$��� NP5s�gN�;Pl�a��%D�d��*Lb����Al��P (&D�@�!.3V���'��@�=I5�$D�t�!̘�L��PoΩB�h���#D�D3��U:vr``݊Rt*� �/&D��E�"/x�1�W�	"�)$%D���iҾ[?��EM�0���D.D�4��K��dlÍ^�=�`� �0D�\�u+Ak���(��^�6�8�+��*D�h��/H�>� ua�"��e�)D��k!�厼�u	�xR}Q'D�$�0"� RFABr��	}@�9!L7D�`��S�-���0��&g�j�*6D�X(��d�.-Hrg\BppR�5D�Q�
�U�$�J�,Y��.�bE(4D�h����*LD~M+�� '���s�6D���!�0��4:�)V�z��$I5D�$���U�C �x��� DB���%D��b6�H:mA�'עDڄZ��!D�� Rq�I��~�Dc��
�)�z]r�"O*��-�*$d�c"��[� T�""O��AQ�Y��9�fe]�g�(��"Oh!3tŒU"�)�T�B2"OFe�i@<6A@q�ķ!�ta&"O6y�ԥ�s� �A��8t�"O�	���ޠ�%F�:2�ܹB"O\�r��J�����&G�32��8b"OH���gκjT̔���$4��hg"O�	��� \^ Hpbe;����C"O��"C��Z�[U�AMՙ��.D�|��FY\�u�`oټ=D����,D���[�[�Z49d��( �!��b=D��	 J
/��U
�N,\�lw�5D���5ӷG�tЩ
C�����"5D��;��Z '�-�t��7s�f����&D��"T��=�l���KXHl�W�$D�4�0��`�m�S�Ӳv���.D��+'�Q�U���Y*<��`)D��ȴ(Z
6�D�e���aPu'D�����[Z�Ѓ�Ž��(�3D�<j���\�������Y����'�/D���b�n����/Үz���H ,D��[妌	�8���jQ"º��(D�� jR9��R
�/8���d&D�8鄊�8fU2��+Pu;D��.D�����Z�T��ٖ�~�L��@�,D����ȣn�����M͍dq��d*D�h��/Ԟ��Q�H�yf���E�&D���R��n
b*��D�B��Ei��$D�䩔*Lv�4�r(��Pp�؉2�#D������1��Q�ԍZ|3N�BR6D��2c@�j�t%����8V*��H�4D�8���\<,�ժ.-�����(D�����U)Z��� �6H�V�ȃ+D� ��>e�DPNA�#r�ad'D����AK@o52�]�������/D�l�DF�h<  �̀(X��@+��9D�`dEQ�'���"��A�Д#uL7D�ܚ�jˑ|��)i1��c˦pː7D� y"o]I�٘�I��yq���e/5D����&�U9*��E��3�4��B�1D�0�͓I	l*��W#/�(���#D�l�q��a�V���S#�h:P!!D��Y���J �����}5E��-:D��xCNZ �Ĳ���Ϥt�ȓc��)ɧ��4K�t�����I�j��ȓ<V��(�D�8"��q��I����&�!�$
�R���q��+x/�T�ȓ�F���x��C��&6���ȓ �Y��JV�*�G�#i?�=���X$A�I� >�yg\�Y�P�ʓB)�eK@�C�C��lk��^ #2�C�	�"4��J0C!uX)R�H�C��C�	Q���Q�	�J��4�B"�[��B�"v��q@TH%�xxt�D-��C�	#�N��˦	L`BG�!sC�C���C��Fd����l �=�C�ɦK���Q��9��١1�\cApC��$U��ǃ�o���T�u�TC�8XVY� S5C7�M�N7n�6C��sv��@F/Pl�	�l�RB�B�	��,�#ED�YzY�1��^��B�I�{�m��HL1�Nǹ6�B�)� z��a�?N@��(TJ��(�|���"OĘ{�T7x��̀`��J���3c"O.5�N�	�����פ=T8 ��"O^ɒ��>KȚa*�C;&j(��"O�Qe����U���\-|�`(�"OP�x�^Z��mA�#����q�"O�8��cCL|:����9��94"OXu�Ҫ���l�0��"5|��"O:��5�ën>�����:R�H�0$"O*,!�D
y��D�˅$���ZV"O�	�3�ٴ=��x�*��� z""Ox�Z��t��|���u�XI!"O�-�ad¾P�4|��(V�:�2,#"O	Q��ʾYd�5�.%��9��"O�����L,J��_ m�R�"O��A���%���*�O�7x��*�"OXh#M�L�ZBIږt\��%"OrᩇO��W��cs�B5<yn�X"Oxa��ُ[
�T3� ��2�d���"O�D
b
�X0�l0FZ�m�ȑ(�"O�4�b��:̜T 3�K7<��Q
�"O�]17ꂁG�) � � E�2�Y�"O����@�u`��%�L�U� �E"O �b(R������(���"OPI���.E}�t�����"O�C�e*ZI�9���\H��DR�"O�ͱ@8�"8(�G�j�S"O.4r�=�	����l��
�"O:y���=s���EԽA���`�"O`�;� Z�qi�Ve�Gk���"Opp�)
�g�0�j�#�?5M���"O��C.��fmB(��W�QA���"Ol���   �P   �
  �  N  #  p,  �5  �;  B  iH  �P  |X  �^  0e  tk  �q  �w  =~  ��  ׊   `� u�	����Zv)C�'ll\�0bOz+��D:�DLVbneќ'�6��	�x
���?T��j�!�45fd��/���I�+��M�TP7��:X�X�i���V�#S���� 7��pLQ�.OM"r�d�>jܺ�ᤨ�8x��lK3I� �u�2-��u��$"A�ﺳ�-���7dI4$��6+vq�(�n::�":j����'<�OLl����V��Nӈ����'���'���'i�����ΉZf� ��4��X�W�''��'���'4���'��y�e_�D��u����F@�7G<cO�&Ud��	ԟ�pc�]��F4��<yoW�H��7m}��T�'Qn,@��L0\�.U˧L$���a�'f�*�!���y��!-6j-*�%���"�@tl�f�r�)�L	=��t���r?�O��n��%��4�窥>ivB����}����5�)�B�v�	�����؟t�s�,��p�$�'��i��N�3} �
s��C������'��7��ঽ[۴n����'���ɤ�s�\�m�M�]�v��b�
pp@un&�a s�IY>I"�oE��v�K�c�/mלГG��Y����H-<Y�K;w��ʁ�X�p����?qA��Ѭ1�N�+�%��F�d8�AJ�?X�D��PBܣ"qT�J�A�"cU�l�ɖԔbC��L�Xl��J<X��i!AM�0T
ɺ��8Cƨ�6��Lkjr�,@ v1�0	�I�����ij�@�-�8�dI�Ӣ���
T��AӢShΙA�a�G�V��E�!e����d�[�*Ԏ 8IMzDP[w���q�X�
v�p�A��Ć80P.i�E'3a��%"#^n�4K��ͪ$� ��A�!31!PE�>0�E�\wĄ��(͎D!T��B�9ɲU���\Y�j$��n J��̋��.�b��1j�T
Di������G��`�A�G��̩���Z���:b���p�W,z�+O��`�(��'@�A�<qY�)���'`�x��M/P��p��<@Vd���	1ZǠ1#%��w�	�	�꜃�d�2	G�T:�O�*����d��Yi��'��	��^q����*�<�� !Q�A3��d�O��D!�)�'}���� �'f?(Qp6K�0�-�=A��~�U���;#��iT�� *�`��,�2i�*�
�޸'�~��6�0���~ͻ- F�#rjB!V���+��I:0$��2��41ˀ���9��q�C+&E��0�u��/�!򤉁Lf�Q!�ؠ-�@�b� �-��'�ўb?݋uh�:.��|KէY������<D��Ђ,	�j
ny �!(����D9�i���
�(O�D��E	�!����A/5��죓Ɖ�{�j��y�	�����nV��B�rU�M�ČK:=���I+�	F�~R)U�^>�����B=D���FE1n�Yz�h�N��:;��o��(��I^"<*�ɩ́�;b �J��.D�|k�oR��&M�&e��B5�<Q�K�7n#����HO�c�\����0pm"�+1�\)�����On� �č m�1Ot�(_x�[!���Һ9C/��S����kY�n��C�I�wvRL)���F��	�Q3A�~B�	�FfQJ�(\'���d ��=Ŷ@�ʓN `�k$�#`��rî��'���I$��'N�B�� $oL�T�#$|mX�{B.�IH!*6M���� '3�tٳ����t�8����'�<���>I�)�7@�ۦ$�H\`�{ӏ¦}��W(V�
�����KУ D�a�4KT J銣<9Hյ0�\e�Ս�+7"�m�'�P��1ct�Y�j��EȖ̘�" ʍ*���q�t�<	�i	��d��4OG��'�Ɩ�5��$�z��cs(A��?y���?���?�M~�yb��� 
"��"�\�d��EH�M�͸'/�#=�Odr�9�]7%�N$�B'x��@�%���b�W�w ������ɽ��n�'Y��L��I�#Mj�|cu�ǀF��'�8�r�ܶ�p<�ecW8L`A�T�W�*� t˘p�<����0A{Ѐ�5�# N� 0!�A�I@���O��<�Q�hx� �H�w9� 	�'�8�K����&��p�ɪ,li��^i}�L2�r"�B�&�+��c䄍"�PP)l������ȋ���)��!���P���<�0-�	�@����F~��U��J�	�Z�#��+}��	�0=i�.�j��BuZ�+{ҩC&�p�
2=��IM�v��ă�nL:����^�:Vt�$6?	��ٟ��|��؟���-)πa�eiJ-|��"� Z�L%��O�ѫ���oMj�
�(��Fl#@Id�, �K(��?!����ۦb���s�U�J~X��(L�u@�;*BON�tr!�i��ѦOL!c�N1�x��'�AL��MH+�[�!�D�*)���5�Z�f����O=��U3�O�{riT�"�1f�
Ӱ����(_b2�O�(���!]��P��LȶsXЋ��'����� �>�$yقl�v�
HX�F3�����Onax�D<�~��'M�	�҆�����s��Łbe@��'}B�i�&|C'o�O�擎I�#���S�? �)7��_�D�U�ܽU�����'I�H�_���'AR�r!�6vYv�3#e6��	��|H�����	͟,Q��{:�J��R:���
�bNy2�')�OQ>��&H��7BMPp��&QuxR�8�ɬ�HO�Sm"����i^�8��Dؓ�ezf���'��)*V��	�y�'��9n��	�G�J�KE$�GKh=����6H����aFb[T9�԰��ҽv�����?�@d�Fhv��7Hֈ�1�<6�M!��<&M �:�ؚ�U�Z%~���Ol�O7���@�==iV�I�G:��y{�Oܠ���'�7�M�O��䡔|������f�S��7P!��NhKN|�A��8� ����Va+Q����'�����dI���թBQZ� *^D$ ���On�d�O&A	3�Z�e���D�O��d�O�A��c�̸��+D�2���T�$�]��,i{ �'.�)�CS<]�	��1O>!fLٷpw#���Fy���%�
[�P�j40ODt'� b1�1O��zS-ł,>� �턙ɶ ��h�z��' �T����j����'�Z`�î��n�ԙ�$Vb����"O�ٖ�&w��2��Hy��J,�y�(��O��u��O�;i^����>��@�'&��Qi��*�B'�<���?a���򤏌@�z��}>���'B�X��0C̒�;E�)����V��$�ꋢP�����4LO�rFc>?*0Mj� ߳$���!mK�,0f] ���o4�*�'�(��U*q��HՄ�6H�lp�5�^��?�%�iY�6-2�I��Oi��s�	�F�U��E�f��)
�dqO�4q���~Ir��׎,�r��G�|⠊�,�����/�}R�O#�[$bU�����b!h6-J*Op����?�1O�ma��]'!!��3�-v�,�A��3>!��J�'Sz]�)�s��[u��F9ay2�5c��;G \._���8��
%�hB�I�U����6h.+�|)���	�HhD➤���?U9��f��L"������p��8-qQ�@�Q���'#=@�O�J,�pJA8[���h�yK �
N>�d2y��U��c�hI�6,\� 7"�����>4�C�I/ude�5eڲ} ���C�/��Oģ=�~��n���F͝�Z��p�@o�<��M�v��@���@�[VL�;��n�'v��"�Q���(����(
^A��1��Y�.r]ze�d�&>��[wF� �#���R?Z8�Tߗ���ѥ.��Px���"O)��p�M�}RP���iZ��y��(!����a�B�+p�ԫ��'�z��(gj���-,Nc�HK' W��y����Q������;������_r�,��'gT#=�T�$U���̠�a��e���a��*���.��C�y�ǒ�Z��!'�	#a��d���`��X�'0�ц�g���#�G1j�J��K-[&!�ēy"\<80lǁ� \��J/T��$Q"O���wIH�d�H {�CĿp�NPc�'1&��P�/l�@;)���(�`2�3�HO~t�T�]v?�$ͯ&%XMе�(f\6e@N�_y��FϦ�h��D\1f.q���;G��P,�i��)gIs+�"�y"���,�<|#��A�EpX\:�K��ְ<1��A�_����M)8�T}ƈ�z!��ɤ��1ؑ
��n��H󦆒�qO�aFzʟ��Ǡ5Δ��������g���(Ox����_�wr��'<g��'D�!��q�E	3+��I$��R�3[/d��dC�[��s ��L�혐� !����D����:#�2���U�%׉'�ўb?%��fݧ{��mc��1?+p��e-D�( �˄�\(թ���+|?��S��/ʓm��	�(OX`zd �����g��?hd�s�A��M��y�O������*~��*�e^9h��!�Q"~\�T�'�h�����sd
A��j˺(t2�'舲�I*4g|�2�͍u �ъ}b�'I��A����W#��C�$��;{�D��'�툵,�*
��I�G�!<��� �r}��3ғ`�qO4�[u&��8m�8+��F�wp�I ��'��(�"�U��'����#鋲��'g��1���5FH�Ƭ����ʆ"O� �BP��D�~��ƪ�
>��
O����X D��D`�ĩ3An��Qf�v�<�0�߽V��2nй@���!Dp��t�{b
V��̹�U�h�F�*�0~[qO��FzB�.?a�I�M� ��%/�BF��P�	�<���F)E��u̓*����}�!`U.�󑦐��X�s��Z�<�g%^�w��A�W���P �xR*B}X�TDyR�]}i������C�C��yܐ�X�h񡁣P
�Ps��ظ'݌#=�Oz���C+4��<aB�>#]�u�6h�}�'} xq/<�I*z�ӫ;����� �d6�I�N
�u��O�Q��A�&K�x�%R�A�^Q��r��4�b��yR(�<E����ۼl1hAf���ē�hO��v���gս~B��
 賒"O���#�^�}���k�g��;�bL{��	���D�O�'_��a�O�F�l9S�G�Xi����ʘcy��<i�j[�OB\�mN�D��6���|��B������S
O��1��n���u��X@�j�"O�dEo�3/�0�D�۸J:�H����,\O
� �
�l���&8�-��"O�)�h� E�  JD%Ę�ա߾���]l�' n������{N��R�5�ވ�K�Oɺ!T�1O"��w +11O�����َ��5>���G�(D� [vD�A�l+�"-F�h��G�&$�x���;��WԞ;����a��1�bB�ɕW�� 2d2PE�%ѤJ�"�Z��$
mܓ1�L��!eW�v&��;��1$���=���I(&�:ms�'Bu����!K�&��e�K� (O"��I(I�1O�Tc�钮u����؄Ȗ8����L�!��ʏ&fl��N_9��Pi1BË�ay�IB/�л�&�.6١EG2Q�6B��7<�������y1phc�Hۅ}8�\؋��?%"�E��U����[�| �X��Ρ$�Q��I��C��'��1�O�%!�+��ɉ6ڥ:&�Y0I>y��E�:�^����Ij�)���ã#nP�%m�0�JB��7�y�&�&d�F�iF�dl*O��=�~��Ѓ��oB�RbH(s��h�<��F�9%$� � ��:f�0W� p�'��j�Q��J�M\�R�2a����3"]��s�H�:XТ��(�b$�I���q3�&-�$l����7<,k�
O�ڷ�G(T{
�����54ل"Ox][��Ѐ��AAD�L%��`#��d7\O��bB��!%�(���"V�\5`%"O����H�m�e
r� ?�ܡ�
	����o�'�|���Q/�LI�=�`�9�o�O��#G)K�^O1O��k�)��"�1O"@2g�E�i5:�#�g[�N.�Ц,*D��:��ȡ=�f��5"ǒ'U�#$$��1�l��Ew��5h\�~��9Z$�J2�y� бYH��YD��~ ���Ҩ��p=��$\`���`��o�V�q�	�}�qO�=yqѬi��ȟYƒ�@g'H��!�ÅN�m��'�zL��1�I&Xp��>�Cr�@�T�]�d%XT�`���-D�$��I �@�&��S2N����,,OD�<Q��+J��؛��W�i�$�c��Q�<Y�&��@��$[�(X���-��FPܓ,6���'K��x孜?�pՋ��.ݲ���n(ʓ&�x�������	 k�Y���!��݋�퇳^��'NHx�-�p<��mS> �<q!������3E��e�<�K��z�^��F2,����r&Ad�	u���O�l��cB��eЬ=v��J�'�)9U��11���@�8�*]����]}2�0ʓ^�^��JT3;���r���Fpd��&��OW�b�<�� &s�VjM�i�03�&�V>�ճ�AQfQ4���$�-iU�B�RBLa�-0�����S�? �mHֈ\��U���a}XF�$\O�}��R�wh�����%�<�{�"O�]�A\�`Rv��rB�5��M��c���dQk�'zp��wHU*Ld�Ay�L*CT�% �O�O�`���+811O�`1$�CJ�1OTa����J~��H��P�Q@�i�"5D��#C�F�t����,g�4����2$�<���P�Ffi{�X!Ŵ1#��yBK���ha�cB�!�6a�!cׄ�p=a��15-��0�	,~��jW`�@qO�Gzr��>���I	6P��kޥo� ���]Cy@�}��� �Kh�n\�}�	�
Ew�D
�o�<a�D�+��m�<�fmɟTk��� B-����nX��Dyҋ���[%hG�~/�E�Ձ1�yR�<ɰ)�#��H�.�	�+����'�|#=�O!��Ʌ���D�"�h՟i�6�cIM�'��(3rA/�I�H�����FҍyU䐞Zv"�c8Cr>�O����lE�.��x��5]\�‍�>u�j���y".��r����@L�g�T�%j��ē�hO����C�CK�v4����8�@=��"Ox{B�ȹl92$+	��D"����$�I�'0^d�`C���̒%�[�Y��c�uɚ=�<��-A�O�1oZ�	����JMd	J���4|�B��G
Od@�b�w�8�+,�Nw"O"��Ț�Y⸽@��J3$��i`�D4\O�E��キ��[	Q5�dѠp"On�I`�FU>	(a�'Zt@�3�F2���u�'�O�$����zq\,P�ƶ�����'�R�y�(���'�^�I��D�Ƙ'������U�݃V�H�@�`��u"O��� &�8Cp��B)A��J,��OA!mO � �P2iL#\�(�KR�<i�B�c*(	h��¡��-J��P��X��{���Cr9.���Q���#�p��=Q&�	�S�py9�'jqy�Zi�l����&"���(Om��'���1O�����	9L ���T�CވcJ�>�!�d��l$�����<�p�����G�ay��	�1��e��O*r�����b-C�I7k�(�7�[5l��i
�h+8���Ћ��?����Kw���B��D�آX��::�Q�h�C`����'l��P�O�8� �/���]z�Lŉ98�A�H>���ٿ9G8 ��	2��ժ���0=����#M���B�	�#���Eݍ!9T�x����B��O��=�~z���a8@��o٧B(��8)At�<���Ǆ~��h��
;3hBH5�Xh�'�n��Q�T'�"�j8�`�����) &P�"ݙ�$
&>�!����zSC���s������69��	�@;���ƪ���is``�&�V���� D��#����^lBS��{<R���*9�I|��ؚ'�ҕo𸊂H�.P�8�:��)D��1�ҩs���H7M�6MXÇ�
_0����HO���=�Cb��H��2F�30��cS˟�s��^��c��{�J�!b6b�H��i6RU���Z�RA�`�E�<� �Ւ?��`��ߡ-����i�uH<��V�$W����/H3
!�r���4�!��ڲ@�MY�郂U.,��"�[�xF�z�O+��"�~xs�P�n	"��Ue���l�<E{r���`�	84$����<��Y��Æ��ʓ'h���s�_�@M�}2F�
^�TU�7��9|��e]�<%�M*t���z�j<M�P,� DO]X�Fy�L�2T�Yb�W�sg������y��3y�TA��8oze"e���'}�"=�O�`�{a�Jx���g�6>[�}ʔ�Tq�'0t��*�I=0 ���Rt`�9'
J G��%GR	*v�O��سJ�g��xRFG,D��mY0kI�R5�I�$\�y�]d�i�����Lp4q��l��ē�hO��� 9R눴!>�Ȩ@*��U��*Q"Oؠ��ɗ��8�5C���h��ɽ��DSz�'�>5��FM,�< QKT=�:4@dɍ"�*9�<Ƀ��^�Oy�mZ�F7B�eM�()̳��+��0��
O�4j�	R�n2�ѣu/	3#��e��"O<��U��-: n@J�ml������$%\O�XwC .�xG�Is{����"O���V��$�H�x��~�aI�K���ğ}�''��x闫���/�z�XT��Q�P��
*=X����O��b�yR�U!1{)���݀W'n� �ĩy!��Ūn&zt��ϸ�����M6O�!�Ā	H� ���8Q0��I�ϖ>���ȓYQ�X�'�7Trq��� rm��I���'��"��A>Fm�T!�оtX��{B�I#z �K�'JQ;Z�4<|2S�H(-����O<��d� *��'��#�����W�����A&0wr؈b����y�`�ј9����,j�h��ÕȰ<����ˏz��<b�� -e���/B�r!�d]&R�����0p^�4�1ctqOx�Fzʟ�Ta�N$=|Ȫ�&5�Vi�9�(O�0�c�g�d��X*����F���j/a��$��`ud�o�f��?nH��4 QQ.�腀�9!���9����Q�0V�8AV��7@��'tўb?-�!Dֲ"94�m�,� �(D��!�K�O�=,�=��ّ�&�e����(O>��d
��hИ��@kڼF�S L�^}��y2�̧�����t��8w���W�F�o���ŞU��t�0
OL(��JJ:;zBh�w�Y�q2`xt"O$��N	U����KP:��-ٗ��:\O�貰aԛc͈�PaT�E�tɑV"O,"��b�bU��Fq�p�y������Xb�'@c����M6r��!s��Z�j`K��%`r&���P.����'�vԑL	DI�9�6o�z�B�w'��z'��A�~uRB��8#�ܹ���'kY ���R$��'�BAۤ-
(.��:P�`}��Y�z��]�;#���e"�	3p����ě�k,	J���zҐ�%>-��O� #����D�֯`y��@�=�f�J��ӟ�|�q�C�u�Ta�ϕ$n�fQ�BBzy��'.|u��m۝5/�ع�/�$9pI�HB��T?��w'����∆4	�@����1|���q	�<��Y�J��'��O^څ�I� :�X�|���g�J�h��av����Y�%�rt�G�ڷ���O�ܔ`de׶���t�*R �,F0�{�l�?VP6�8q�p�c枤'���v}���Olr�|��%_ZP���	Ga������'��)��6?ɳ�ρW�HR���/&$	13��~�<	��(�l�{��C�^3��`�/a�a�d�� ����Z�*x��d#[Ă��x",�	��H���'b(�#�G�Ɵ4�	ȟ��ɰzn.( ��C7f�����#�A`���i�~� ��OY<R�)�� �)������JB�����	Q|�iM�o�Yq�םN&89���F�$ b@w��]�6�?#<�%��-�$��\��3��C~�kX�<����hO0��3#����!�M6EiE�V��.RB�	:�,Q�A�*@�.Uڶ��-0��x3�'�,Q���OqT�d�<Qp���r0��
&���	%��xG: ���i���'��'���l H"=�(���K8�pE	��? �2,q��a��L��[4��d���.<O\��c@v�e��ʖ���sР-H�0;��Y���a*҆���<��؟�{d��2halcr��,��5�!ʟ���s���h�^� `Л6�Ab�f=6�J�;g%O�Gy�oU/�ܘR��!$ʌARD����U"���ĺ<�@�JW+>=�'�?1�O��ܣ���"߲x��/Ǧ�H!��OAp��̟��	l&
�	6H��\y�X�t��xݛ��	��0�ל	}DR�d_:~B̀��D�m^L��g��eN\Tj�V�t��:iN4{Pnޜ�Vك,C���O�P�1�'k��	ͱvh���%��[JвV�Y"��ݟ@��ɣOe(l�ƪŮL����pI@,H&�'hL"=�O���	�'r¡�c!O�̶��V+�0�9-O|�����T��D�OF�'D,���?��\�+D�����Z,�������?I���0{&�Ҷ+Q<L�X��?%��gS�n�x�O� �e��-^d����j��%��'&����x�|��%��>E�d��{\����`�.6�p����F�y�%N��?�������4��� �I�.˺k��%��H����"Ol����1S�~�9��M�'����q���<A�d�t����,�7y�@	�K�?U��P�o� ��h��|2�y����ɿ�i[g�C�����X.s��I��<D�L�D�Ɛ � `��%k�y�E�5D�\ȕ-��z��l�!'�9k$��X��%�$$�O ���ȧ;ކ@���UW
 �
OX�y��JF����4.@��&�3�~o/ғ>Q��J�BA��A7�F57�9���ֹ��$"<��%���D�+7����@Y 9���;p�h1D���v�Ł=-@�ha��b�d�1�O��	�!
 ������4T����)*��B��92�����@J09-�2��Y����d]|�'5�t�d#$���@����X�0H�В�yҨ�/J ��0�'j5�
9�W/^C!N��5�ϸyO��"��'�
吧���y)��'����dk� ^+�L��I#󂭫1��/T'4�ca$� k�#>YV�Si�O36ب"dG�e(�a��гd_�D[���ƇQ?U	�㋐Ka�(pA�j݈�j*D�����oI��&DrT��%�3}
#�S�T��&�~(V-��;F��aU4l��LϾ���O�7��f�|�i��?�d�z���c��0�%&��Jwp|[�yҁ�S���O� {�4TH4�q�� �ѫ�Ƙ+>��aRQ%�:M�����F,b��ʣh[�Q����+�p��qV?e�;v�̭aա�O�����:ܵCg��AP�����ᦑ�I�v��у�?~�^%�I֟��S�?��@��l�G��n@F1c�옧4\���
צ�M���O̐]�FT'�y��%������ 	� R����daڶ��M{,��*�)fl�a�V��?A��K���k��S;N����O�����\�	f��9`��h�@�E'^�`����#W���OD�"��� 7��Ik���s�����
�J�88D��n��i�7���P�C&2�'��m�4M�"�)�O��D���)G�5��K�8 ��"$Kڏ-��z�nK������O��"�P�{�'� ���M�;��DH`vP{U��aw��H��T)@��牷R�����OH�R�^L��)�O`�����U8��4fJ�3���gy ܀�&��@���Ͳ6 ����O�`�;�ʞ'Y��	��M{��fŒ���6b'�`��.綅C@fǁ�yR��	�?q��`l� �V�����?�B&��W8QB�ԉsE
Qp -tƛF���?IxX�eȢ
R�'w���O��ݫZ���J�H�!a%�O�)E(�@�.@	Du�7MJ�#�"��PN�<A���?�����=��P�kϘ��+C������S�<�s� pl⃳���T@�G��' "P�|8��j��O<�ġ�P9��0BGTy2Cߺb��"Ģ>!����D�<�J~
�'�>�cF�%������5=ε�}r�)��S2k�K>Q�\��29�=�	�'W�T`uAԽCi�s�a2Z\�i	�'���B�Z�u^�i+��)]y�[
�'�͢�Cѭ4[���IQ>P��]h�'�d0��N�(L�2Y���E��	�'El�D��3�%���i�n<��NC�<��m��B� Yr��h��+c�F@�<��
�Dx��P��鰔gINy�<q��@��y���L3_jR�ʳ�Tw�<)A���F��80v�]0�x�{��q�<�c'�h��Z�&�]b�XR�<�ph��M��n��@�$iVF��H�"���Ж#�@C�ݲu(��* 8=��&R�����¹��p���-7d9���v\�k��Ia��� ǘ<f�x<���ϧ �F���7l���i�S'�qsȈ�g���F$�N@�5��9��H�vaA$N��K�
	cE�MX.�Si�'��A鍵tWQ9��@U��4(
�'�z���;}� )X�
��>�n�3	�'%"H�W�П�)��9(	�'����{�P��h�d�*�'�ڄ($A�)$��ݡ� �]��
�'$�Y�JҡT�4�Sf���݊�'""��ş�| ��Iֶxf�@�'� a��Ϫn0*U�"�R4p�e#�'~�B��%T���h+|A��'���f*L�s������;_l���'�f����ܖ}��pd��"jɛ�'0�tʠ���0�r�J�'�m�H��' ���GC��:���^�2��q���� ��c�?���Z©.Y�8��"O�(q��2O������OS��P�"Ofi�)�7&�ڥ�姘�@����"OlL�Q���Pi�2W`��2b�W"O��� B˝h��1�o66A>�qw"O���/ֹ{�������"L���"Of�#��]&\I&/ڍ*��@��"O����܅|�:�a�-/{���U"O`�悌  ��e�J�"j�"O�@����s�`1��AtWNH
�"O���g�*�H h�`�$ZtHE"O��
V����j��DE�� "O|!q0�݁zk���3eT#"u��*�"O�ye`�%zD�� ゎ�.rx%��"O���pi�"W?tXd(� a�4��"OB8�e	��hH�f��"o�d�1C"O^�)�Ó;7�0	1�в6��4�'"O��B)�)\�J���.��3�RP#b"O��BJ�;J�3 `��v��բ�"O����"k��Hυ��Չ�"Oօ�3��Wޔ��3�;u��f"Of�
u���[��EK��Ly|!qt"O���O�e��I���GKT8xA"O��h�Ù,�hё�B�2'���y"ꎝc�����<Bd��1��y�T�kU�(�#�P�_����Cf�D�<	�m��d���P��R�8NH�䥎o�<R�R#C2��U'��H��D�W�<qvӭ/��PB���=Ș`�D _V�<�w)�jm��9"�	�� �p�V�<4* *g��e�p\�#N�y7��R�<I4��&�ܑ;Q���5媩(R-P�<I#��F�҂f�QT���h�<a-��=��ܛ�a�.*�����e�<I�Rc״�F �3�0�)�iBg�<�2oã`�T����ɞA��(S�`L_�<Q��c!$p���$Mw���%^�<��kZ�z�$���!�L$�r�-�\�<)�l(�.{�hQv_r*�W�<��P��L9��߬$�2�i�#�S�<��.d��A�6���&\�ACJ�<�q��y�z�@"�ќ>4��c��E�<�G�^�`ɤ�0D�E255���C�<	a,�!�r��� �	C������B�<�q,�"y�x�㤏 A�H<����}�<�cNVu�B�!���UѴ����}�<iCC(Nt|`��M�>�:Гp@B�<I�	��p�lI�f�J�'xa��{�<i��;Ğ4p��X�"X�$$�z�<aw�_^�="&�!���n�]�<aS��0?�6�8C��FA@�cl�O�<�dl��8�,I��횯D(��RR ]q�<��7d�L���FK
�JnOj�<�G�Mh�YX�+�	,~+�OXd�<�+:��PZ2���1���VIE�<i0�K"�j ��^����Ԋ�C�<���� �p�v�˻B�` �,�Z�<yW$�35U�y"(��I�Ҩp瀚K�<��EΑ^��%Jm��ܼc�LL�<	��G�*�@����0(���� �S�<���i�X�g@X�I��PiS�<�SMT g0��b��FQ���amVP�<ѶD���n���ߡsh��Y�CJ�<��&hX2��UH�&	�6�Q`EJ�<� X5ʑ�ʒ'CD�oԢPdB��g"O�ؘ�'�8�8�p��0*O���"O��aq*ف��� �Q/0:��ڇ"Or��(�VC<"��[�Q. I{"O�d�* �0t$�9�Q�N��І"Oֱz��M7xR� b����M����*O�MY�N�<;bL�0�|4	�'���P�D��0��<c���9�'#����<6TJ�sI[�N���'��2�%�M�\�-�����'ʐ�h@�ϟ=��z&�)���'�h%ŭ׉dX�<	��ɮ3
�2�'����+�������_0V�Z���'�:q�JƤcO����fݴ���
�'/�!��Oݑ.�V�F�
����
�'����+���%p�-�5F���[�'O04����z�0��ho>J���'���'�zR��є��=8.�,��'`�g9V,(�4���5*�p�'�B�
�F]9;��C�و,v��{�'��c�yq ;6���Rjh�0�'GL����P.A���[�I���'7���Ӣ��(��9���9]� �'(&�#[|Y�� ���,VP��'�v}pql����EnA!(m�1p�'�T� ת�t)�MI��]^]0�'i��i�F�Ծ���h��P��'=XTI�K�i0�-ұ],�Q�'1N���E�NG�iå�	U�΅�'Z��
�-��lc�l��O�$z��s�'ϴiY�E� H�f�# 7�A��'ʄ��/��]/�� �CF���'���#�;,��aPa ؜?oz5z�'��!>;�ģ�57d����'��D!�ˑ)V�4�3�y~�T�'���W�T�H��
�rnА��'�Č6kW�Q��$Z�C[�b@�e�	�'���A�D���C�k'DgR1�	�'*�h* IG�
�uR�O	�95d2�'�H�F�����rvj0$k,U�'��5{RJ7J�
��eG�e$���'Hn�)',(�>��R&JW�u��'CZp�CN2 �ܑ�1_:&��X�'=~m)�ȴr�`��e@�5<܈c�'g��"1/��]��Q��%4�I��'���Q�%�L	�-˵G�$9�`��'�:e"�^�jJn�����h8��'�|����A*�}ٖG׬bU�5�'bBE0%�v��٥CS�q�Ĺ��'F����?َժ�f�$���'�����3;����fA�]/��r�'���ɲ� :�HH�E��AX
�'��LyS�Ԫ��J2��G;X��'���)�JĢG]���/U�	�'j��!�O�:�* Y4l ::Շ�4B={f��c�sGPx�-��-��{q��'y6d�xP�O�6U�ȓ)��dvh >]h���h�lzrхȓX&�)"pЄ��H++X���6� �*D�<^�!����(�N���Mh%���	;�&�����7v.Շȓh:��s��a���ě�g�.��ȓMe�T�CO�.Q�����zn����5���T-ϙK��L�� ��ą�S�? �`�-�-��ɺ���/Tݖa[P"Od	ɰ�0є]+F��>G���"O~p�C�3O���L�/u0�2�"O>�tM֮Z*���K�U�T���"O��I�!�r�z��(W�fEf0D��;��J�xT�3ᐦzK:4
�,D��+�L\.��Ǣ۫;�8��u,D�hzGK�<0�D	q��U-*�ܐ��5D�����	>�p�sv@	���H.D�T#sD_�D���[r�ٖѾ1��)D����
��z�����AE�����"D��S��9P��
�<=xPZa�3D��q�67�<	���,?�����%D�hH���AS}+��)����Ԫ#D��q'�$=�<!󦂹¶�Y�.#D���#�w|p�0"�pz�`g� D�K�@}zdc`�3�$�qD=D�ACF16����'眒b#�9k�<D�(ѱ��-k����GY�x���֦&D���,ɵ���
�.$!�#&8D��i���-�b�
v��+q�8W� D���v�]�,}��g�dݼmY�&?D��a/l�֝��,T&p{���?D�X����!�8�$�d�2p؁k'D�8���9F�(Ua��ހ ���#N'D��YpDK$A��`s�W�Qt��q��%D�����/�����иWJ`<[p�6D�4jj����(d%�B ��cT
B��*������g�au$���C�IM��hCB�
!�p�*1n^O��C�	�m� ��PEe�>C����C�	0�Hi� L�
1��U�lT<C�IG�����L��D�y�T8�B�I�;A�S�Đt7��PՃ5�B�q|�$�
5��8�I�	�B�'*�4hɁ��0
��&e��(��B�+����V�O5:p#m���B�	�F/N��/]�{;Њq-A�RonB�-��{�����y80H@# ;C�Ij:�����b�0���$�B��<��CF�_��\Kv �r	 B䉔T���Ӳń�'Y�t��H��3�B�ɓH2�}CF�غ��D�d͘'J5<C�	�'��a允�U9D���N�
_�C䉐1���.]�� ��^4�%��'~���&�T4q��̃^#D\)2�'.x��CC�M�j�pt�v�ZYa�'*�`�4ZG:51,�%v>���'��3��� ��5hՋ�-��'����� �D�N(@�ʗz�����'W�a(�޽�X�a��}k8Q�'|xf�����	G�B�t����'���D|.ܤ���F�f�1@�'�Pi���?�~�u�p�6I!�'~�<ҢLܙX��a!��-8ot�b�'����f�z�,Я5�Q��'Z� �I�z�\���ԫ��a��{r�ݑw��QѰ��l���*�fO��H|��ISo����u�o��5����X�L"����p�d[��ǨtjB�I�e��9����C�
,�0�C!d��B��	��Q����N
�C��%o�B�I5.�"=s�7Vg���ւB�j��B��<C����P�tU�C�hB�h�n��E��vb@a;�j�%hTB�)� �%҆m^��NM�'�	Ej���"O8|Ӳ�� ��z5[	�����"O�=�W��& ���I��2#"Oz���C�%&z\�󨔷~�X�(5"O�y(c
��)c���%�CHʆq*""O����郧j�B�(w�A/V� "O��œY+���-_�04"O@E��
�Zn� ��+j��R"O��;fE�R$�@R������'�y��9��F�I��(�����y�] X�L9%�L�g��P��y�*�.[1��b�_;.��i�e��$�y�  e�Đq&�3ư�%�݌�y�IO2S.�����Ӏ,̒dn��e�!�dȱ:m0YB��M�Qh"ͪ/�!�Đ=�ʩ�d"�=0+н
d�2"�!����
�2�*�%at��pC�p!���$:�p�D/E*.��=r���!Qs!�=c�&QS%���T��P�o!�$�0{�P�7i�'2y�������rD!�� f`�Zր2;pP�9 N�v�!�d@�\F�xڣLW2j�Ix0��$*�!��ԻYp�Ӗ��8O����6�� }!�Dق@��M�m�z���f�a!��S�V:�h�Ͼ^.X)p�A�lB��i�G��FAz���&���Mk�I ����Z/�z�ہ�ϣ����H:N���Ԧ8��i2'��1"|�qmŧLE�m��6S��R"��:��|�V`�v�',2وʃ= �$��ׅ8,8�qJ� ����Ձ(x\qK�&���`���P@Z�w�[,Rf�J�
�,����&Z�V�[T��������{0��Ė� 
0i�!LE�l:���(�\�b��IB���X�9�!�L�<��a1���<vт ǈ��`$H$ɡ�c��b)��Ms�,�3��d�32�ʜ�A/�L�tl����d���-��h:'�
�%�dy��ɎP�P� ���S�*��UG���	��E�'�����%Fb����
<�1j�f"@����O1k�*�}����pONk���h7e�8����d/,(��2K��B�G.���r���#J��;����'B
S�D�p�*X��	l:���=��ܱ0��H)���d�`q!�D�J	�mx���j���r
�`��᫖dЖ�����B��Mc8��9��$�l�0eOO�V,�I���٭T ��E�JL�Q��W�r\8A��xd�v�\%��5Ac-ϕcPd���Ov�'΀q��8�~li�i�9]�,�sϓ��lh�m�)}��r&�w��HZ�eX E@��pW�S Sr(�r,����'û��a�b蚕FxN}AH���f8�}@L�{=���ë�	�.Yl:�iQc181Ka�(O�ft�����<�!�$�ML��#vIW��<���N�d|�ƀ�,B��%Z#�ۨ�Mk��$����K*3+r�CE�#��� �H2k:��d��rgNy����Z0��e&ޢ<~�)u✇~_g�8y&b-�Q�N�'�~��B�S�	��09�B�%�ϓ)�"08�F�T������ČږAx�D##X��)��-�o���#�D��*dɒ�J��	I�g���j�4	H�c�|rA�B@��b֬�o:�i�4��#�%��8��E��&^�!��x\	P  !�6X�s�Z�
�pPab�υ E�0�i���MkW�?�ӽ��+���X�GJ�CмI�0l!@O�I2���-c�$	)R�0������$c���3�H��u�) ���!H��IG҆�>>>5�d�G2+�����<�f �9�*���q-(袓G��A��������I!�N�G94���'-f`��a���Dj���`x�*L>i���@8j+�f�)_�Py��G������5n���	�_ڂycB���y��	�%Jx�\-N�����R3�0�R����H���n�Yc��Py�-
CŒ�I���+Nw�)��D���xb,F�f�{�Y-S� y�CE>l(�`6l��wA�3	ȀWz��&'� �\��@!p���U��S� ��ȓ{.�0��&I-�茋�b¬<�BA��S�? `	�W̐��)ѡ�A���0""O�� h��M�����d��P��t�W"O�x%LU*pd~�*��2���"Oz��/\���(�kP�l�u"O����y/j]3d*�N4fE	�"O�%�C�~D�p��P�zfH1"O(���MP�~�Y�O Z阕�Q"O���-	> ]l��ڽ"�Hd�"O����ʰ�F����/��taP"OV���CZFl9b��X����"O� ׃�* y2�m�,F+|�RD2D����ڿc,��bW$
&wy^�P�5D� [�"UC��9C��L� �R�2D�찁��x�Lty�H,Qd$���C?D�HK�I67�l��H7E�� C�� D�$	w��>�����$f�,�-.D�����Ɏ5�܍��J�5Od���/D��p�#��j�RLv��!&h��9��0D��PG-6m�y����]�:ѫ<D�Ȫ�'�7$p'AO��={�<D�D�%D�R�&I�qG�:�%���-D�h�E���{	bh�T�0iV�a᧊.D��*���'m��i������q��*D��0�؈w����ČU��B���+D���5�+`�������j0����&D��`'�-P�h��J�V�[��%D�P��"=����B
�V8�J��.D��;5���b�D�yT,��'k��2D���ݱ):�)����3>�H1%0D� :'�	�4ތ�%a��&Xi��>D�d�A[de|�2ӆl���>D�8�����]�#��w/����<���&7���􄙈2�@��ߍv���B�ߟ��~�&��q8�K�2ML4{ o0xOJM��Ӵc9!�$@>�:\2�`�IZ0H1�`��l2ў�
�߁NL0Z N�v�'g��`4/Ч_2]I��X�T���ȓ}V�T7�;hG.����`��I�1ʱ�r�҉{A̱�����5(�-/@p�]�Rh�����*D��RG�A**��%���92�!C�h�?��M2,+�!�(	��3�Hin�c4��#wڽ��I_�J%ta��I=�*�ҁB�`��q�FC�z�8a#+�[�P܉�i�>'�4E���	�^��� R�[�H-�`k�6%�T"<ѢL��E����CCQ�p7��Xt�&���^6i���p�QFB!��ђ�yRa/��A2���w����H�'t�Fq���Z8d#j�x`��< 4x@��9O�xXլ��J�f�E���\`p"Of����ΒOЍ���F#/C�kcn��x��-���(�l5�6쎑vf����+TL����;�(� �:����R/@n.�i����=E�N)5Z<iAN��Oܐ�޳��P�5�O渋�
����{�-ĕfR����\
���s�_���#�K�k���'-K1 Bi���j%+�G��S��E�ȓ+��jv���^�
v�ɱ&o���FF^�&G:`x�䕈 ��i�.	[�O���J p�zl�E���E;f�dq!򄘢;� �(I��vԚl[c�^9Z�(��
�2�jC�ٖuFQ�O.���NA� ���I�� W`�dJ�D*�O� '-Cd����h��l9�7��a����dkȒq@h4ǆ��p?��g/�D\ӱ��H|Ј�t�]^�'n��G/�$�T���k� ����z�ǩ��a�ኀO�'3�rIG"O~�"t#����1O\��10$\�z� �9b��jp�1?E�$B��ak�tOE�"M �y"M�B�:Qr��ϗ-f.dz2��Rtʓ~߶����ٸ*x���'��3�h6�hр
n�8G��W�����m�:!�­@�J�}lH���b	h��$#�*D(!���-m L[�ǛYKXM���S�b/� s���)��y�%c9�Sg����� _r����ŃU(B�)� ��׋A�)�`ɀ���*G���p��OL�C�f�V�O�>��$1�2����	�!AНc/D� :�e��L)>���X����a��-��H�Q.���*Q�6�Y��==�:"tm�5xb!�ğ�jrr!8Wo�X��6����B�	:]���ڧ��v=$9�2LK\ehC�ɴ�ԑJ`e�!d�R+1�Wze4C�	
Ҫ�@��3g�4#�K��b�C��j�Z �B��R��#���/�C�I�0�����M�*\;��t�W8Q<�C�I�����Ѐ�As$����q �C�8o3h����m��5 ��tC�I�R0N5�㜬��x%�ŅPgjC䉊�H����= H���q�B�e�\��bA<P����ɀ�>�4B�*J@9d���n����@g��o�B�	[�0�sG�.s���R�̟��B䉝F� KB�]�*�H��ю�S�B�	�6�a��'у"(U��C�K��B�	�=�
@��W;Rߨ�Ԥ_�C��B�ɕ.	�� ��$j����[�U~rC�I� )z���PP�&-���*5�C�ɗ8�a���p�$}�6	V�yC�	*4,���1+�� I��C�	y&�U1�cO�XG�q��lΟ�B��(F���a�>A�8D����h��B�j8����?w�L1�b�#,��B�	&T鴨�	ܖ��+�#�>t�B�I>`���E�Q��#�EfZC�	�0<�HXqA]�Z����BMI�6�LC�	�)��}ӡ�A	/;l1*�jAJ�(C��3Z04��6+N��bR:>��B�	�̐���:a��%Z�Q�fB�	�%��p�,DՒ�9�8��C�	�C����_�R��Q�����C�	�X��ȸU�ӷw�J\X�^I'�C䉳S3R�8�*~��b��u��C��#|QRɹ2nS'tT�UQ��Y���B䉫VT�չq�I5�X���w�B�I8{�y�〜�0�{e��L}�C�	�	�2嘗oK*6�0Ҵ
h�B�	#Qt6�3e��_��u�ԺNrC䉬����d\��TR!i�c/vC�ɫ>|�E�O	+f���ǵ<\�B䉶m�
���5fR�8��D�*�B�IE�xѺB��'�R=[���`�.B�I�P�$�uj���LE���H��C�ɃPk0�{%GNz��	1���m+|C�ɵ7 ���g��S�[�rFC��7�<���d����doXd��C��H��I���2���t�7Y<�C�I#<N����.��Ah�(�o�C�I�C�ڥ@�!*C���R���3RD�C�I�m�*L�|Ȍ�0�͸0ŠC�IJ@�d[&���-\-�
�1)�B䉪���G���K��C7��-j�lB�	2S~��&�ُ�z��_�IC�I92����#�-
�`G�S�)}�C�%!��G��(@�M���N���C�Ɍ;�^��p'��N���t��K�xB��8��m@v`I:5�h�
1]l�:➄��&F]����j�#R�D�>�d]�5�ʹ�T/U7<B�	��J,j�!�EY�����Ɂ�w�ι㢮G �!�dN,y�\mx�C&lj0�Kd��# �!�� \e�S�_�	�p�`c��Q{�('"O�l�����;����iz��X��"O"�ЊE| -�J���q"O�=hՁ�..I��AWj����"Oj��#kĨ}J�Ո�+b]�]��"OT�����&�:�y ��%9y@M�C"O6����8r��kDFĨUtʐ��"O�b���b�<����Mb d( "OT�g�H-v��m�d�'	.}!�$Z0L� q�c�gSd5�'/!򤕤>x��RP���6r�1Sw�˜B!�D�7\:l�EfޥMa����-�h�!�Ěi^�k�%YiT�Hv�G��!�$�MĈ�%�6/Q�@$�ѧ1�!�DJ�,j�K�"եb;�ͩT��3�!�$D�"�(D8Ee�T) ���=&�!�̙T�H��=�H(	Յ6u!�ĖGz�IS��
2v���W��6wc!�$��@�L�	t�G<G	�&ǘ�d=!�U�!��IpB�\�u�ĤIS�֔Q5!�dѭ91j�WlF;c��$�/��3�!��^�	צ\���BpXRL��b%!�d� s��D"PT�URx�r�k�s�!�K�d!�`���C�x�'$�UQ!�M�����T(T>�T�hY/7T!�d\�"�P@A�V6Z��b���_�!�R\��#��KE��s�;�!��ҙ2��\x���Py�4�+O!�D�4񦼊e+X�O�v��U���!�dI"X���V�X��KEĐ�We!���.�I�����A5)�␢~y!�Ċ-D��DĪ`Iu���2T!�D������NF�����ݫ>B!�;o��㇍۪b��-��ެ_(!��#29^U�T��#hxܭR���	�!�d�!�P�R�m�BԠ��D�M9R�!�$@*-_�����.9Ǧ|�%�C&�!��@�`�(}�0�D!L���#S�!���u��M�"�� �Լ脣�%=!�A:i��2���V�����S!!�ğ��H��G��G��	#�#7(!��2$�ȭ�"Þ2=61P�c��b!�@ւ�
�Z�2�A�-{!� �=����.^�p�[�O2b!�Րw���@0l��E��8p���|�!�䁁J02�W�W9G��k"��K)!�"b��Q�d
->�i3�gON�!��������蔙��R��!�DB$y��� �,o�|�� F�H�!�$Ź-�l� �9�"�m�b�!��P7*}F���Td8'��)`�"x��'�l%AA䟙Z1�1�aÆ�#~�*H<i�k�2H��B�FjF��'2��ȓ�`YX��
A��5cW�K�4�U�ȓ3c�
���K�6��Q�/>Ƥ��k|�sn�3g0y@I��X�1��'v��;g�JT���w%²wn�#�'N��kWˀ�Mv�(WC�tj��'b�p+��B�H��/�1x�ȥ��'�|��AB����fLL+:H�	�'�.��N��d����E�'bVps	�'Sz��QE�Q�$�����.m��h��'�̨0J����I��`b5B�'K�U`���q�"�� ��ZHJ�"��� 0H2�� ����8N<͈�"OʬS��u^�L�nѤ)Tjtq�"O�-���S�OL����?�<�s"OU�r��a�P��S!�n0��1"O��13`��V���$�`�"O~������"(k�l�*<D"�"Ot]��+ă[��!�3�!��i�r"O⵸�Y��m�3ږq�v��"Ot(�@ՐXUYf$�*t��a2"Oz b5���W��iv�H2d+��{�"O�x(E�,q�����j�vA����"O���f�_+��`���+*�A9�"O�t�6G�> ��3�%�n1Г"O:p�k�&��	YwD�F��I!"O2EK�[/J3���b�W�|5�"O��񅓼77�Y��C�&rP��"O���S �E���AB�mb�<�W"O��[�/P	<~� ҥ6S>Fh�"O�t��� ��)y�b70ܩ�A"O�I��дQ�a0�g]0�	�"O�0�4#WF$� f�2[�>�2"O,�r�̋�K�e����jŰL �"O>�k�kע��=�!&�����"OD�Qd�zP;�嚥9�-�4"OΤ�a�:��-P�I��l��"O� 3r'��R�A�$��y�"O��QW/��j���Pe�!�"O��0cT�}����aa��̕�v"O �7)�$a���;�`٪orRA��"OFH�3) #t~�;T�U4m�	�"O��Cr���r�x��Q�P�_�HI2�"O�DSd���f����"G�;C���I�"O6u	�C�����[��̌����"O�t��>>�^4��"�Ɖ�7"On�tE*DK
�䄟`x0a+"O��rm� ��E�i]���"O,� EکDQv�	E]��d���"O�Y�ͬ,�2E���	C��i�"O\p�J�n6�0�I�Dr��"O(�`'H!h�;����(���"O��0� EZ�Ƽ���D�y(�"O,l�gjۧ*�L	2��3��PT"O���bH.~��9{�[ /�`�"O����.g|��w����p��"Ope@$ב90fP�&��h�xd@�"O���sӃ0	�ʤ�^�*qȐr�"OtY���������fr��A�"O�X�����%���H���ZwDU�Q"O����,Ux���"O�FF
�Q�m6D�t��,��V$�a�L̛3V��1��1D�|��ёg�r���JV���K#D��8�a��ѫ�.�+Q�j}�3�"D�L�����74<QZ�B�L��Ц#D�\j���7m�´D�D)欪RO!D�(��%B�.��Pxgԋ])�xj��?D��Y�cA�h�.��P�_f����-)D� ���m#��b��H'm�Й�<D�4z��� J��pH*x�7D������0N6p�׍B�f�
� #�5D���V�4(�L`�(��#��4D�Щ�L�#|���NǑM��Q`�2D�k&� An��MF:{�j�7�.D�tPq㝍� 1�q�2�R�y�o2D������.>�Q�l���X��1D�� �A���9`���
��l8��"O04Y!�W�� ۴l� ��	1W"Ob��f�d-n�1Ū�/�8��"O��� J�5V�"�y�\+i�e�"O����l��z���y%j�2x-L|+�"O�`(�L]�Et�;e�L,��
e"O�x B)J�sX�b���b|��c"O uH�Θ{ڌ�:��:��,V"O
� �B� Q�LR�&W�:�`Y�#"O̘���yU�eS YҜdY�"O�XB�H�V�D8Ѓ�,Y�<)bd"O����hʁP�HE��Q�S&9k�"O�<��b����K��'4`i�`"O&	1vi^�&�nTb�*�m&p�"O�D���&2����9(Zu�Q"O�A����=�,�8'��;R"F�R�"OH��� Ԟ)����u�Q=Mɣ"Ota�ƅW�,�&������"O�W�ЭN��|a�-X.j���e"O��K��ߣ7¾%1PMػd1i� "OT��G�4WkV ��FӧxM$	��"Ob!�Z�HҢ� a��i���)�"O|5�B�F��qQꙶ&�j��%"Oi�Ɗ���	)a-`ђ��"O&�%�ꬌ�C�P���q"ORL3��C�D-����� z�g"O��{t�Ǫ5�d	A�)�CB�"Oz ��k^�m�u���[70��B�"O��)�g�CBޡz���2o��"O��1W�I���/[&��7"O�i8�K�Dp�2rH�6GHt�C�"OH���儻� iKG J��	�"O
��#/�u�d���F
A�h�a"Oꔓ�ᘙbܹ[�k�	6 �W"OjE�#h`Ɉ�;6����q"Ob�ْ$��8�}tMƮ�^�1t"O�;%��u��˔�B��r�kC"O�p�gN%4�b� ��Ng�6�b�"O�@1EX%t�����C�{��m�g"O ;��@�/�P�@s��&��(@�"Ot��B�ilNdKĤ��D\�"OЀ��� �]r����I}�8�Q�"OP陓k�Y�vT@��7ی��t"O�� `����t�t�Ǳk�<�"O��Z��Kv�\�H4
Z=~�5I�"O�i���.9������3x*6"O�1��.B��r�q�玍V)�A�"O��uƁ�<���5}l�1B�"O0�cgC�D�$U�3�+b�:7"Ox�'i��T�j�%��t��"O¡�C�^EL�(�$Ղ�`	jc"Obl�#l]%9-^���MR����"O֨��扭E�V8C$�'(�!��"O��3"/�%I� :�"À[��A"O:s�.E���M����#M�R�XE"OzlCĂ�-�j��CP/|o`�a�"Oܔ�Po�/7��[�D�:}Hp%ل"O��
cŀ-�FP�D��9����"O�us��ʅO]>Q�� ����!)�"OFu90m�}?�53� �$�R���"O�=+s'�P���h�d'su^-2�"O�I;T�{PN���un:��!"O<��Fʃ1��5)�kE3^���"O�Y��<ya�Y9VE�6e�dbs"O� ��0G�Vg�@$1��	IQ`��"O`�k���S��SCͬ?n��Z�"O�e)6/I5Iu�)C5��Y\�H�&"O�- �oǶ',��W.kJu	�"O�`��f_�|d��vmJ� ��"O8	1$BM{x�d�7=F��"O�LiWeHg�z%���	�w)ʹۢ"O�C�@::l��o
4p"�"O��D�I%w7R�yu�}Wƀ�c"O�ي@l��r�n��ңZ*w?܍��"O��ZGd��p�����>r�� �*OV0�!/[�2��@{��C�+\fb	�'�����D��V�φ�@iA�'�H}�S��o�#tE���P���'��qA�I��(^���$�:JI��'�����L6+��qpD�ͱ-�a��'a��`��`$��`��	Rhc�'h�P�FO(��0��i�LQ�'p��A-]�M��"́f{$��'�l��DcH/&(  m�>}x�'m���Ǣ@�_��eS�ȥ~����'
%q�a�*=>%{���|Մ�z�'U�y�7��0hh�(@�i�&sP⥋�'CbX����fj�)AhK%l���'�~��RM�=^�Y�+��k�h�'6ƍ�C�\mXQ���^� �k�'�6��ˈ$~���۬ ��1R�'�,)k׫�)�X���ޔE~���'��K��ˬe<��!�I˅ �\�;	�'�p�J�U�#2 ��S-	���*
�'�������x�Ԗݶ�
�'��1%*յxx`a�f�#��
�'V�|���@6*Vh���b҅gػ	�'������
N<<L�p�UR�չ	�'H���"�x�@�)���*C�B�+�'�t�6-�=@h��FN<
`�5�
�'F�p�$�©1����AM�L�:
�'U����9R<��A�> ^YK�'�^����ċ���!�ɓ>1����'6`IA�$S�A��&-����'�Ȥ�gNJQ�4M+���4�	�'`�*$(D��
�{�U@h��	�'̠P�$�G9'�����Q8<�|`�'*P$ÒB'(�8Z0	W�׮U��'r���d��G�8�P`m �x�t���'b`rwF
�B��\�����_И�8�'� 5��RjqiWB��"��ԁ�'6�[��{���bW�Tc�<E��'#bM
��Ԗ'�<Hz��YZ��'+�X����.fLLa�gJ<K��8�	�'�>�5��#4%�`r4-�F����	�'x�����C֝�d�/']m��'�L@��]�E],�S�/�H�'*�h!��q
���(�.ܰ�'2T�vŏ#�$�xe�Af�)�"O��IRJ�"\n�bCJX�C�X"OF���+I�~\����) >'G.��t"OM@�D�b�Vy��K8d'�9c"O.(1�D�Ox̔�p�I>{�"O�x���t��DaS;z�Bc"O����,ŋ8_�)'a_>$�A"OhP�7�ɭ%O*aТo�4[:zs"Ozx+���k����o�>7Ө���"O�x;A��\C�����"�n�R�"O� b�ذK��,ox��D��XϺ��"O��K�V$�F]��.,�=��"OZ�`CI����5�+�4�6"O`Q�v'� *�=�#�B���!"OH	0C��;u *��K`.�"O<��G��Q�䙃�o^)�v�9$"O��*�ϼ)M�����|��"O<��0"���P9��̺�����yB��j�m�@�O�(���yr�@,F<%S�(A�8eơ&I
��y"��#w&�I0��=7A>(�I&�y��>c̄�@�#Ǌyi��y򌉑E>$��+��i,D��y��m���󦙖=X���
��yr��a֦-x��N�^X�!�4	��y���(�5kr�I0T@I�Q<�y���XL�9�sLY91MCB�V.�y2��J�ؑ�/߇=���1.�)�yb'�yZZ-P��ǥARJH"r��>�y��G=h����I�8���I�#���yү�/f�����#��P#L�ybmC�7���J�';F�6xSS��#�y�Ư,�����/_8kz�2��yRI�^�м8TKH�Y�2��cK��yB��!1�H�r�R��rd&�
�yR�W�k�9�R."���Q�y�c�; �̽0��8yq>�+�,�yB��$}����*�xǞ0j5A��yb��:l���uK	e�ԝ�D�W>�yr��!@��y�
�\�|������y��@�m���re�<V����UH�	�yA�*gP��BFY2N"�k�ܹ�y®��w����xK\�PU��y�o�,7�It�\<:}������y�EG�hq��"{��S��W�y舴4w50�o"�����	�yR+�&7�n%
��٣�̀�`���y)�.d�:�L�6	��1�)ߕ�yB`��+��t8���0 ����j�#�y��B���%u�nx�S!ˌ��y2hO'���&�S�̀N��y�G+tj�T�r�� H�21�-@+�y�삹��):����B{��z��y�D�'0F�@p��9�@�H��[��y"�Ô�tir�M��/ܜd�q@��y".E1x��@钪!�� �/���y�Ռ	;�ɷ
R�1T^�8���y��Xд��B�#��H�Gב�y��Q��(�D�:��YWlҚ�yRL�wd�2�b��Zx��� �%�y��l��q����:�r�y��A*�yBeY"j)�Ļ�˛��u8����yB��1f�iZ�*�0	d8�1���!�yR���h%YD�ր�>,�a'D �y�凬PZ��<g34\ ��?{�C�I����p���-A;�	cg�.�.B�I~<�Qe�<-��E�wR;�B䉏d����3jό-��lB4U$6C�"	�1R��V����ā�H�FC�Ʌ<�T8��ٰw�"L�@B�8PTC�I<n��CK�|Z�C����|B��'�6�2���"���d�]�ujPB��?K�����I;� ��%�52�DB�	�qG���ϰ�]p׈�IBB�)� (�*��
7DL����^-s(���"O�ܨ��@�%A���*�)��A�"O�
6D�<�LAY ��c����G"OِE
e����C<aF8��"O��S`��g�D�1���H��"O��J`.��j�����=D
	3"O�0���\Av�8U����Q��"O��S$���m!3��/'6̸�%"O�
��R
�R�e��.�q��"O�� gZ$�$�
�I�y�Q"O�e�i�!8�)�IC�԰ v"Ozs��W�Aun��M��ẅl;Q"O����']�BV�4�Wٛ)��ܺ"O$Ђ4��5���
�%�Հ�"O�eS�3�(���	r����"O��p��Ϡ3�\cď�=�f���"O��������A���e~q��"O�Y�ԇPjklh�Ǫ�gN�z�"O�tscS�b�!��Ș)���"O���C�(P���A�fA#� ��"O�=�rj�:S���+�$)��I0d"O�a
���;2�ꀐ�J�M�\iе"O��SC"+^Ͷ�Ih\ p��$"O(�%�=\�b��G��j�LA�"O@�Pc)�*�Ѵ�V�IP\�A"O��C �؄ �ċ�55P�q�"OB4����yG
����ܘ,@!�$R8GG��J�IҶgE��7ke%!��Ʉ,�9�V�L�v8�D#DJI=�!�׳C̅�BkS�ʞ�`f�>�!�$�V�4�&�2F����D��.�!���&����bB�*�j�0����!�D@	C�,�I�'z��� ���\�!��ˌ/&��B��NT��l�u(��%%!�O��2��ӥ���(=f!��2>%ɣ��. �^�y�!�!�D�>zx@1�R+x�@�.3�!�V`��E��6F�>m�a�в8m!�SA�,ٓ��U<([��
0��	P!�� �f)�&T� ��0��d!�]�p-8$���^�>��b̓�!���V�4b'Z�i'$|���R�!�d(��,�bg�0j!�S�!�$��;�Ai�X d�Yt��1�!�$��i�8VN �]�jM!��!�!�$ߧ}�b0�m�<� ���f���!��Q+��3��9-�:-THǏ,�!�D�j��B�!�FԺ�K���<�!���Y��@6�	�"�܉��Bd�!�_�;���1/�4�u)$��n{!�]Q��0BF-�Y�~C�@�.�!򄌗3�$��F��Q�l�#�\�G�!��<d��t��h[$���P�!���`wx�٦Z/R��X�C���!�_�s�)+��܈�L�A�/�O�!��B�mi�!�(��@���Z�!��Ȉq��4i0�/	{d�։O/�!��Ψ0�m 𥅫)Ӡ=���J=#�!�..�ȡ��������`F�z�!�ßK�P=H�M��)?�I�Jl!�	�ɸ̐��
�%ƴ! �Z�5�!����p� 7��
v������e�!��s�TXpi�:8Բ &�e�!�$�9��8�,Z�Tf�=Ӓ����!�� j��4�#uB\X'��:��w"O@��u`K#
�p��04q��"O��٣��}��퀱!Ϙv�l�"e"O0�`6iQ0��r'a;A�]yt"OH��bÏ�q�ǠĀ0������⟘j@�
��؈��K��|�8I�w��//�Q!2̍�M����^�������&ىe,�"|�	�,v�}D@�p�D[0MH0��#=a&	I���9�Y˓��dH�$	Pp��_�5�����HO�T���'725�)`ӴS�%
�&�CwC�}Fdܑ�LK��?!���w ��b0M��JV�P�B?�0	�-O��Fz�����ЦMmZ
sa��j�E9�|5���Q�R�.�I�O�6��%�I�T���)�2��'�ddS�)~ �x�3K�j�l�M��=Q�M$o��	����%ғusf�ڑ@�s���)��k��<moN��h��@������v���T1rө�2&�<%2����MӑA������M��ň���U->����Q�(0TC����~��'�ўl�>YR�8)�R�kvd�=B`�@#��`�	�y�g�]�(7m;��O���]�(V@
��<}R-��L]�I�B-O�4�7 �ͦE�?qÃ�����I��L��I�[��]0���;�d���(��)�mѬ��C�&M����q�R�x�:O���W�:
������P���$ˑQS֝�A͏�[�P 2(�2sQ�Ik��$�OR�'�8��ş��'�5�$M�bv���v��.���!<�S�O����P>Ow,@�B�FD�<Mb���~Z
8����M�K>�S��*O��i�l�%L��i���,d�4d�>׼���(8��2n�2c�h`�l�I�UBpс3���:'0|i�o�
Rz��SaW�jȡ`�/�O�� plL�Ѧ�f|x��˓)a6�-�sa�A���8B�ˍ�<Q�ek�'4����M3�`��X����&�����Tas_�6M�O�ʓ�?9�*�P�e��&Dn&D2��T�d�2��%�h�ZY;�M�rV|��V�.�����\���M(O p� �P��;���'9S�Ta1�d�:�N�����"��i}�����<��Y�	h5�Tw��?Y�)Ŕ}'�T�K3���5Dh�'i���e�ƶ"f����5��UQ�y�Q8_n�2�" �{�*#=At	����	���'�M�'nƊAc��zP�߷!�`ZR9x�f,�����|�	�I;�9Qdˑ�����D$�pɖ��<��~��A�N��i�V0��w�$|Q&(��!�>��'6B,8gኄ�y�R���8W;V�%�<� �
�t���qBn

<Z��RPe�3	j�����''xϓ�?�'XX"<)����'|�ٚP �� .��+c�S�!;�bC b3�Qg�/Jd�����i����I�=�J�SEČ1(��l۴2~�D�I柘8�4�?1���i��BE��9Z V7�ǮwM��a�Oz�d7|O6ۣX�pɁ<��R����
N�'` �I�F�	A��L8nZ�1z��#�i��h����EO�&��H>Q�[t��  @�?