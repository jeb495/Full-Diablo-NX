MPQ    ��	    h�  h                                                                                 ��I=H!
ʜ�i����n�����t��3���;�D��W�>S �5�!ݮBv�"��ݞ�r<tB��'�r�����zٝ�0C�?#���Yy���*�>�wȈ�i/��nt)xWOo�A�3"��o_����V�N#}A3r�ܥB����-��8���[A���S�*i!�lH��_=L�;�����RH��8 MІ"�����C q���������蠖�S�X�y|�p��'�+��R��4Kx�V��⸔A� ]���bq�Yu<z'Dvm�7&%s
��b�� %N��!M��	k�!N�It5�X�����05n��0pHD�]_��.n���<x)�	d�At�+v:�5��ħ��9N�oC��*�_�bN:����z�~���Qs�T|�!*�0s�L��F��* �{R1׾�I�`|n���<����Q-��p������Oٚ!�����f��B�����)��)���� �#�X�R��]�f���[�^ז��n�n����8�SO_��Vl0~��"���9CܖV�ɯ!~��z9tI�Mr���/�/՚��ʛE)�Z<�V^Q�Ђ����!5Ҥ'�5bනd^,���\sQ����+T����W�V�_d���y����n�=��I��`L�*VJ	+�b�儤}L����si��^!����5X�l/Zꨖ�@���Q��q6��.�S�9����aG_�V9.13Il�D�Ģ<\F�|]yE��$Ӛ"	�~:�:�|�@�o*dSK����}XRT�0B8�2B�!�o}4��N���(
,�ئR�/ha١�u�7N ��0D���c�y��)Q�4mCܫ�wm��#�#�T1J5GC��#��r���0�:~�
��޽�G�Y?d�h����>�~YoM@Cu�����<ގ��<t,���t_�)�VqE}Y����� {���8	,� �d��̙JkU�n�L����	<1�-�-1���@j�x�K0Vh��-�!��:,�Ŵ��IV���:L����`3b��נ�iؠ�8�E��2�������HZ�"*����ٸ��O�yx�m��(	��1�O��P�.���c�c��&��������7��$�7�T���Б�������X�1�G��z�"ϽlR��'���"a��,��/��7�E?��C��s��n�8������E;/ӗ]50f���]�"��5�~P��G���Z7�\{+8Z�F�r0p��!���i˃��/ҿQ�S5bhj9�jq��i�f��s\F7t�Ŀ>�d�V�qo5�>��o|�N�ԟyVTY�ƌd��H�4h{2�rJ[%�~|M7�[D����lh��@W��B�������D�Ġ�]C�8��x$�Z뚫�GB����T�� ��{x.`�aM�	}�:�&w
��"���d|�W��3���u7/@�џLc��x�͓��i*�x>������*�P6�������8�ga�,�9Ʉ��*t��9��U�&��Q��'��ȓ
<���/�Ղ��Z\P����H��� 4��&�sA	�P�4)�j}�fi�C(P�-�<p�����R�E�a\��ޏ�3sч-�"y�����ou]�}F@ʏ*^㇣2K�Jr��M��j�}���g�(�Q��60=>�� rRIs��H���T�E�ܒY�4��i��C ���lH���^;���0�VR���H�ߊn)�cN
B��� ��Z]�h�BUdJn��. Q�~
:��Զ؛ K�<D����v@��X�����o���t���.�lp�jok���ē���g1���U�@�����xo�z��-�h��z��V�2��U���Ϳ�#k�2MNC�،Fmu�o]f��g~��wn�D5F�Bw�(Z!z�I�7�d�
k�U�G��x؎�P��yR��+�}���ڋ�.ʲ�ƴe�ȿ��эW�0?&NY
d�.߼�]�>O�dqxҍ	���T�2gJ�tC4gݬ�C�k��V�pP¿(�J*���|n�y5a����o�Q��`I��\�/�,�`ݣ<5��2
��I���e�X9��uI�N�
ҿwL�e�?^(�CWGjmH(�� ޑXy�?��QSx�`���ީ��v��8�s����{4���{����l7���޶�!��=E3̳�^����D�$��穃��	�B�O� ��)�ܡ�'
W�
X)y|�8e���L�N;��FՃn,S�[ݯ�����q,Dp���2&�r�e�����y�F9����pr��w�˒ ���د��O�b��=-e����N���؉&�G��>�a[Ts���Ԇ��Xē� �V����I�e�|�(z����B�p�N����F$��а�q��.ϊ߬.=�Q��ܫ��>05f��d��;���+3��|���^�us�!�k��^"v���(1��Zy�Tz��R^�j�mf�4ӭ��B={���EY�˓`�f�b��>���#�7�h>�֕l�
�hE�Xgh67�Nt�(��J��N^n�C^��,wԻ*��B`G��"��wZ̯S�z��Wܔ`��86�6:������`�̘8�G��Ů,�p|^���67?K8zJ�LUET��I&�)zY�l�u�/|5$��4�� \H�OT�+���z��83*���K��xʠa�<�pA۽����)�H�z���������i$��,|�M��1�F�M�H�܈h��=%��&�4�i'�qsf��R��1�Q��k�ꮖ�suL9G�HR0 �4�^r� x�!�c�&��������]RTml��ѥ_	�h)%��M����dr�H\������E�A��*D�k�b�m�d�^¶�uv�bfy k;��hT|6!;A�K�k(� �R\�r��^�&,�2�]����ju�s����<���Z��5��)���M�۳%�L�i���I���ǚ�]<M����28���#v���_TГZC��o��Ccn�ð��RW�����	�-�]��d���beEz�Kd�?ng�?*�Fi�	w����pV�xr�	%�N�5D�д��N�����-Knʹw*�F@������m&^��m� o��Ov�<I�:-)Ry5��]�Ƈ��mcg�xP+p(H��:J����٘��2����&4YR�]�׀ϰL�ӷO�k���\��´`ZR61Ri?�օI�A~����*D��l��!_ؘ*;�t���Hzi h�"&�U��X�q)��d"�����,^EXy�jˋǙ'"���-i�4�:����"�.�Af�]K�m�}��ps�D�37��-.�bn�% Ԑn��{�UPU��c�I�XX_�=��<�n3F0+?��x-#���ΰ�dd_�d������]�5U3��¦&´*����d��y�����:��Y�5Й��ҍx��/��!=�0��u�G�F��嗤{m��9n��;>j�I�;<+4�Le���Ng4��󚜷����$K�窸��$��rП�?�>Hm����]j~d��n��Q>��<��,�qSj�V�ѿ#~��7�"�(�����
�g�>Ztd�r������j������@�C�>���k���r
5��-�p���QmT^'�k����pdh+o�I�q��Vi#w�-<���n�7$�Q<����~L�&AJ���b�T������v�sdp1¹�D���^X�SvZes���ݩ+�����6��ή�6�B�|w_lQ.�cl+�l�=�;F��)y��9���k$&��"�@�:���|�7o�6K�2@�`�+X�&0]�=2��s�J�����%�f�'չ���.h��ې��7����إD1���Zx�f�Q�@m��^�����	���Tl�Gެ2#�kr�Q0�:"�z
wQ��cUYz��h�s�沐5~� "@��۳�+)��E�i]�?��t��)�o|�)V�E8����Uқ��꺪,ҭv�p!���FJ�<)�����}℩���18g�@WG�F�Vår�	A��O7�@m�$�T��L��D�[�T��z����������̈́�@�l�'��C�5"����P;���ߺ��Qms�_	��L��Ŗ�d.�Z���a�c��������S�r�S$q��O�/�+P���x��	��ӆJ���ܵ��XC����3�K��dA~��ǀ�lgE�]U��=�� �n������bo;4�0�د@f��;���;�Q��~K؆���6�b\��\Z�|r�7�32����I���p��p��h���j�"8a����9ȟ�YF2U"�U��դqHUo�y�>���|�tJ�:g�VO���!MΥo�4+�V2+��J6������m[?Kd���h��@r�jBt�C��Ȋ�۠8!!��ζN��x߿Z�ćG�~w`YLT�0a�+��.[�pa�Y}�'r�*�
c/�"iuKdG�3W��3��͂Уk@z�igR�K�n��iee�x���!쎅��P�Kz�ӘxV��B.�,:���$CoS�97ʹU;4��l���W���<�+M/l���Z�6<.��cO��焥��AS��P�z �ev�fĜ(�ϛW��g���-���`�\%�{ފ�n�-��t��������1{^��6�2i2��t����h���;�)}��>I(3�y�1�>>*J -	s��_�� ����4.�ض�hm�l��'�הΥ��:.�1�)� ���%�Q��R�
������r�u���)�U?o��Fz� ��~��Z�#�V�KZa�_��v��#$�?d���]���ݨ l�	j�z���&��΢>��蓂���3���RPx��z���-��c�L{�ج�V�Nvz���D#���g��Nj���Y��W�f�O��D$�2 �DP	B�Zߜ����p��}bka�����x���P�w�RK��*F�Z��u�;.�/@�����o
��p-Ww��&)+d�;]�x?>J�qy�э��  Z"�2B�JtB[gx̝C�~N��[P}}�(̆B*�W��yp��F��/p�v�`:�wcR/����;�9<Uc���'`���I8e^,�����Ɋ�
�=4L�5?���>ˆj�;E(o`v ��|�r���RQ���`W!ޤ��v��8N]����2#�V�n�g�lҺQ���!��/= �#�ΰ}�Av����$�G��K1���QB��r i�T�-�,ڢ�@��2)��y8 !����N\����u������yfC�H�9Dd��-�6�Ϳ��܌��z��|F��nP�������ˍQ����j�!�j@��z�te�1��������&�g>���[����q��ǖ��g�L�`����Ѥ� �[b|���zI6�Y(ԉ(�ǫB'�A��<,ðt_����8�ZI�=�}��S,�پ�f�E��aU��[�3�ao�>�R^�L��\���X�v�����K���T��R�:�j��l�o���L��{��W�s<3��v$`���bBlv�]�U���>�ȕ��:���D*`�Gg~�;6��t�����ӰNY�D�j������,��*q"�B;ʤ�]��w�q�S��	��T)`���8Q��:2���`I���1�ӴI��	����p7ms��?��pU#rL�9@�>Ł&�4YY;�u��
�I��ր�\SG�O�:�+���z� 8�W���0*���S��a�F<p�,��ty�&N�H������2y}柤$6��|���HY1P�NMs�ܣ�ڸ�V�x�p4Q��'_��a�wRH�Y�Q#����)�>�N��9?r6H����/̫^ͫ_ 3�Γ~ ~�m35�����_Tj���V�	O9�%M�1��XG�h��#�yW�/�&��<�*��!�����1uQ���i ��c��6|a���<DkCݠ�ͨ��M�ԙ�P,yM��X�
�U�4�.jÌո� V�ּ`�d���x� �����WQP��Ք�A@�M\Q���g�&�@v�y�3	�N��C��5q\n��ϬWbM�4��.�d���ǃd���bཡz���z���)ۋ�7�d���8pq��rY�s%o���p�	�O))N�����4��~��d�w�$�F�$��F�r.W^����{�`�
5p<'�[:�oaRT�ɔ�4{��жc ����mp�T�H�JJyUY��Y���q��'�&/Á���􀊅���?�O[#��s\�dv��[}6,��i�uȅL�\�|x,�*l�d�_s;����J��H5T �4]"�p}լ� qdf	��;��^����X4E�˦�'��p�Ik4�^��'[��9A�hG]�+�-��O���o�D�7\`� ��b�w: ����жK�י�I���X�����h�n^�0�Ul����$�F΋��[�d%)����3`5�]����/'7��fV"�My���:P����E�д]���w�
�D!x.�0C`�Bz�F=t�Oq{�Lp״ q� v���<��w�G���&o�"w��*d��������_s��E��ߠ��Zh¨Y�I�H$�]E�v��D�콆�*$���a��S��L3~��N�r�o.����e���;"�tr�rn`����̥G3�FEq�;��uA���*�蓼�{5���ѫ�Y��H|^"�����+^�+�,܇��XVDZ�h�$�b�n�Q������]n�L�B�J�I�b�㩤� `�O(5s_U��
�F��X�ZEZ�]j�"��Q��M��6���	6S���3�}_��.�ܮlf%��+�F�R�y��ѕ���$Am�"���:�:|I7o`)�K�x����9Xȕ�0x��28c��%Ӳ��Z���t"斦�h�0�۫T�7D%���Dl<���#��B�QR�jm�I����C�k>�%FT���Gy��#�rjs�0R��=p�
�#����Y��h'��~��@��&�ȟ�����DD�zxitb���j��)��E�*�"0P����<,{W������J!Dl�s~�	J���6��1s?�@�6ξA�V�/�����
�ER����q
L3���VOlC�5�*���h�.�¨�{�_���+�>�"��#�}� ���w�o5�mN�&	9��!�S�ݘV.5d�_c�$��B��|̭��$�J�ن.��~"̈́${V�N����N���Ҿ��9n���,����vѐ��:��E����X��a�n�B�T�eȎ"�;O}�SJ�f��k���h���~F8���I��Ьn\�O)Zv��r�y��nbާ,���n�uF���h�3�jgSx<�W��H�:�/F-K��z
p����� o+�/>`�|���t�VJ�k�|-��* �4F:2��J1����om�D[:�تL��h{\{@�E!B����	��d���7�J��� x������G�B;E�T7�u���b.V�;aq�}����N)
���"D�d�@mW�Y�3��,�+0�@5�7�an=��I�i��&xt?����y��f�P��U������,u*���ҽj��9��U�a.䇩���^�~�i<�/��
/qZ|���~���]��&�A�%&P���`�Uf�A(�$��rƏ����[�	]\��8ޅ��)xN-h��4���e(�������`r��}��2���ȃ�ʶ�}w3g��D(�~¦,�>f�V ���sρ!���H���I��4�迶��6��k�������U��f��[����G��bR
�ʃȒՆ��ᛢ^��U���Zl ���~ ���)��pK4�F�ڠv��	�^��T��՛�nu�c0l�E�j��_���	��)Ö�}Kf����l�6x�Ozv�-�@�ɇ|��G�V܊o�@��C�|#�����N�Z��e���vf	W�+��Dk��Bm��Z�8]���}��|k	3Y���dxN�P�K�R�o�xq�����?b.��3�j��}7Y�0UW�U�&"d"i��>Eumq�&�$8����2d4t}�:gbC������P8[(�*�D��2޽y��p���n�-ў�<1`���Ӓ��/
y���?<����<=����I���e ��,��DY�
�ۀLC�?�	�9_�j#O(*� N�:��aQ� |`�B�ޟEv@S:8	g��Q�*���1���slm)����!ZN7=�<���ʼ%*��6�$�IW���/BBX $��H�?�߶���g)�fX8�MJ���N��[|:��_�QH8�T[&�q{D��#�(�(��eB��gi�< �u\��Wﭮˈ��i��%z"�����Ԩe�|�2��~j���C&6���Z,[9����$��d�	�瓃���o��U<�9�|�djzħ@��������F���<rB��u�/����@���=n��R2�tmZf��1������3��ɏ���^�C���e��/rtv�c|������H�T�k�RT�Wj�����mo��+2{��n��S-�Aya`��b�	�QJ����:�m�v>����K}昀�/{+�g���6�8t-��̀.kNT�J���t���,�l*�UxBm�����w�7QS�Lo��=`[:�8l�f:�x��;� �֡*�n�c�>j��s�p���'#]?A��0�L�M��`$&�'*Y�)Du\���������$\�f
OAA,+���zT&8}��Ʌ��h�.H[a$q�pw���l���)Hl�ջ�d\�#��z��$q�|:���Ct�1��M.ލܾ�.�3���SP�4��'���\#�R���79�-����d�)��9z��H�u��*ң^(qX �A�������e�ͤ���T��8��'�	�)�%����ˮ��������3U�����7��*��w�أ���x�¬7�u,6� ���^!6ק{�wNjk^&��H��(�,��WO,�t�Sڃ�-���Q���V��6���c�䟅%׃B���
Y�F�y���隼B�M7���=-�����v�A;����	LC+����n�����{��5��#d������jd��b[Vzl{�����T4d���ڿ+�TO�p��vr԰�%J��������tN�'��L}��Һ 0�w S'F����XjX��^����5d���<B�	:#��R/g�����-8c��2�.mpp��H�9J���da�!��އ&*M�L�Ez�����O�j	i�\&?��} 6'ܩi�i�����wL���*��;l�I-_��;����ޘH�^> ��D"QՇ�Hq�V\�T3��}Iܖ�ҟX����Ad'����H<4�O�'�k�zVA��]��M�e������UD' r7�-���b$� J�;�2+��K=N����I%	@X�6&�ٴvn���0�����)����9�f�N�w�d��}��K*�5˖���xªC5ڧ]�����S:���������A�҃'��� �!�`�0�®='�F�h[['B{�\�/�֦�!��`<aݛ�B5����� �E!���β�>�������7)�WG:C�V��tr��l6] ��H��/���8T��CDS�������~�����d�
TR��������%(t��r�Lيu6=��]����6����d6�����!U\��`5cOJ��^���D�^���m����w�+�}��gU}V��8��unҋ����hL�~OJz	�bh�$�.�0���sZZ��o�}�(�Xց�Z[h��|H��5O���6���d���]
�+_��.��)l����s�"F���yV���B9�$\j�"zaY:c�|��6o�;�K�����X�f(0��o2�N�� .�:W�QAp�cT�h�����'�7�C�m�AD���4��>�Q��mt0���G����fօT�N�G4�#���r��0�#X�
��[�MY��h��z樔^~j�k@t�U��3�wӛ�K��Z�t�
��e�)�E��{�=��ґB��p�4,HhL5z����tJ|k���M�$�8�z�ȕ�|�1�7@;6�<�=Vy*-^%L�ڥ�6>X��E��tpL�g��Q`s�6����8����Y������]�t�9� ";E��8�������Ðm)J~	t�>�	�����.���O��c5�߿�͎��U���$��J�E���,h�9�d�?|�ɯ`����+KώP������?������\�b&fE����A���D�n|���@��I�;jT���fh���@����,~A�9�X�E͋�\��Z���r�.c���B��n��L'�������=h��.j⣄)�o���Z�F(a��ߘ�K�.�X�o��V>;�|<!M�p�+VE���-"��_4a�%2!iaJ��Ȍ/p_"[5�i���~h6��@���Bj�o��j?���#�n�����W�xU���VXG�WZQ�Tr^�ag\.Q�ba^�}Ga���
Y�z"�d�ҚWQ3�3������@�
����O��$X2i�tx�������;>TPg�U�8��n����'x,���Z�ey9�U���䢮q�.1�Y[�<Sr6/����	ZmF"������"���MA���P�e��[�fz-(��������]�Q���u�Ҹ\[�ހ�8��!-#�X�O|O���ҜG�����x��2\�y�{<Ȟ��1�Y}R�_��I(iEc�'�U>��C � 5s���U����i�C�-4d��|�"p���8��0�0�̪������[�j����
S�u�M𾠫Sע�t;U��ZY "�i~��*���̱KO��U�iv�Ԃ��guǄ��a��ɤX�adl���j���:|i�D��Ġ=�x���Qt�'��x�Hz��-��
�V��^V���f\��3Y#��T]w�N�k7�����*�f(��x1����1D�GB�ݰZ����2_�5�k%e�X��x	ERP�?�RA��Sب������ .�����O�8��0Wm�&�.Fd]����ۆ>@��q/�0�:�=S��P2� Nt��g�k�C���g��P�X�(ы*��FHy�*H�|�2�K�,`z�ӭ��/�-��<����r��y�I�`e�3n�'��G�
c�]L~q�?/��4Zj~��(�}; /�����ЇQ�`UN�ޚĔv��g8Đ׫2���l���Af�l�X��4�!��=v���)��7�����$L\�������B�� �K��c!�ژ����5�)*K86�����NNyZG#��2a�̭~�/p9�!�DA�O�#ǿ���� h;��t����źPη�!D+�H�h˃z�֢��Z�����p��en�X����;�&�=�o�W[T�%��jІZ���D������	�Z���/|�2Vz?9��Ӻ��������7I���x��B�����P��=I5Nٍ�<qf�i"����Ѧb3񉌏4�^�Z���W�ʫ�v�Ѐ�9�oŋ�eT��R��oj^S���jn���{�"�)�G����`2uPb8��,�Ʊ˿���>���֦߃�;�y��~gt�G6ȝ%thc���NOx,� ���M�,�d�*g�6B�/F��مw+S��Тh��`��8�:(����˷�	6�֢�=W�p���BI,?���5$L�4�t�&�V\Y8�u]:�k�U��I\ɥ O�g�+��.z�_�88��t j~�	� a_�.p0����چ��pH'~	��K���U��$�nR|՝��>�1�}M�X'��~�ڮq�.�4�f�'�H�W~�R�Qb=��HC5�XW�e9�(�H#HE�%�w^�V� ��U��0��cj������Y`�T>�����	:�%Ý���^�^�s��M+ʹ�UW��2e�*Un�J����=�'yvu��f <!�Y��62��2�Tky���á����!,�*��N,Y��S���A ����*��'M�,ǳӣ�>�����*4ǚ7e'M��x��\2Cv�)3�����CF ܟ+,Snf���Ͳ�(f���U���Վb�d0�b�GzGCc��WE��^ŋ`h�iY�8p��QrO��%%G���N�Ѕ4�N�pH�吨^F'�w��F��X��C�ܨ^~���1����<]k�:��VR
0a�� �ȇ�c����+3pYH"H,��Jo���?�I�\�{����&%���n5΀ ���w�O�[D�\a9��1�;6"Q-iP~��zk3��n�*Ո�l4O�_�>�;�6ϊ �H��� ��"����bW�q�f��J5�xTh�==�X����ܮu'��"��h]47,���T�POAws]|��ν9�E#���DbFP7�.���b�� ���Mn5���\��e�I`:�X0���� n��0\�$��W��tX�A L�Ud[�F�G��@�5�x�����%�ڂީ�Z_����:��f�/��Ej���,����!0y��8��F��B{�
�ת�Ȧ�C���h<��W�=����}\�\�`�3��<�e��#(�{���-����c���7[�>�;]�����h�ʁE��fڔ�����S�_#�Bz�~_�:������z!��%�I�t��cr�J^�Pb�:�|�x�1y��+�t�BY��<�8����5>�`�!�p�"`t^���l���M+��؇���V�.��޹�UOQn����b�f���2L�rJ��WbCa��i5����psU���r��w�X��{Z֒n�����˸�L.6���ο��s8�O�_�l�.��l܅���*F���y�������$w�
"�!�:>��|���o�nK�d�q�uX>W�0���2.Z��ۨ�u���޿hE���,hM?���7:��H�gD����}Z!Q�!m/7O��%���	A�uT;�G�� #��r ��0ȏOs�{
��q�6w�Y+��h]���F�~�t�@/�h���T�
���q��\gt�T��`��)g�Ei8��XN����K�c,�uU�.���+�Jײ�Z�@�?>����S����1�Ou@�U�7�VԜj�7�#O	�V*��5Z��*Li��L�/�]�:E�՘Ѫ$_��^����������4>`"�M��kx�D��erBm�e	��Wj���`O.��u�
�cP�¿y�x���#(B$B���@�k�<K������Z���D�]�y�V�fQ��)�ꫀ�2�\�i��?$���ݵ1Ewz=�|���߄Fnw̠
���;�Kz�IߺfC���I���"�.~<X}��h��F��\��Zl�r�A��"ۧb��Է��+��?̹h֭-j]]�ԹR�`�p=cF#�T�0�!�'��po!Li>�w|w�����V@�É2N��7�4|42�o�JǼ1�j��7[0O�>�h��@�AB�%H�t�!�0}V�	,�X��_�x%���,G���|aT������.La�a���}.q�{
ԅ�"��Od���W�,"3��^��!@�p���(u�����ci=�x�����i��5�P"�y�S!��n���T,뚃��Q1`<�9H�QUl��������43	<�E�/= � +~Zȓ(m������ӥ�!A�9PSW�V!�fե@(<ϛ�����T0ƾ�1��\����{��ߞ�-ޝ@�jb9�[[��w ,�2�Ic�s��2���69ȹ��ʬ|�}-(��"(,\�"Xk>� ^%�sښ��=ힱ z�~�C4�k����=�}��XGo�;=��Jn���q���*���[����
�I��+��庢TJ�UН���zz ��~��k��؇w�Kjqi����v�L��EVZY��G��$J��ٱl���j] �Wf�媷_�ܓs�g�D>�⅐xۛ�z��-{,����r�}ǳV�b��������#����xN���2�)�(��f�n��W�cu�D�*RBc*!ZpЀ�5����zk�6ͺ�Yx��P�SR�~�._B�h��Fr.�f�� ����&�K=W���&�`zd�#P�I��>;��q�U���)�nq��J�2���t�cgI�C�wg��r;P�v3(��*|����"y!�s�{���'��S`5�/��C�/ �Z���<���r�2�IIۊe�g��Bbo�:V�
>w�L�
�?�j�/��j�Տ(�< J*�D���Q?IG`�yޕcNv�/U8�t�M3� ����̿|Cl���ʞ]!��=1ƭ��Kʲ�G��~$��S�
��`B��H ����~x��4G�v�)e�Q8�q���Nmx��10��t�G3q�
�|���D܊3��������x��y�2�7�+�c�\S����~�,�؛[P��(�����eIrG��,�������&���*R[o�Ʒwё�5	���[��z��ѵ���F�|� jz��7���o�:���|mI�2@n�MO���� �%���Y=$�j����*�f�+o�r������3N���2�^h���j�e�v�]��"�F�=T��RJ�j95� �����{�[qʄ⁈��G`M~b���Dñ�"���d>�ь�ba��M��g��6��bt�5G̶ChNJf�{8�k�,�Լ*��B�?��w�"�S��.��}�`��`8�u�:�����L٘����&��Z�phY��]�#?7���mLA�<��&���Yjf�u�Vx�9h�"�g�W\�Ow� +~�z
��8���2�	 ��E�a�%�p��?���ņ7{�H�A�SH��I�0�i$��1|p���9�91aDEM�����ph�); �	�A4��'0�,R��RY,bc1�c �������9�[H�:�� >(^�[j d�/������5��������?T�"yֽ)	`j�%~���	�����ʴ3\V\����-A7*�o�N�Д�¢�du�7�NWs �IÞT0�6������k�2�>Nl����J��,J��I���fp��_��&���ҢgM��h׹5[�����(M�E�,���8M�"鳧n���(v�1�D���YCaJP���PnA�L��u�Ea�ݩ�u�M�I�dK�CbQ�Kz"+�+;⯊�������u���@�p³r��$% ڔ�!='� ��N����n���6&�w�F�K��<8�C0z^y�9��|K�;1�<xa�:<R���I�чc�c�<��	�p� HG�YJ��iz�����Q�y& �8��>����l�D�O��$<\�SJ�� �6�,i����5+l����3*�r�lot�_D�;�%�[}�Hf�� Ժ"���=�iq�����V�s�����Xef���;O'�-����4rg-�]��F$A�(�]7f���5p��� ��ND���7-)��q�bڸx ��hу�A�w�h�AI��xX�o�Ϭ�no�I0Z��䥷�����A�P�d�sG�|��wx5Az~�.�2 ��]��������#:aT��!�V�jb�yV)��.)!)%F0��3�sFNa*�6�{���%xF�����5��<���8���75LS�ɜ{��V�@�n����7��=���Ћ�㨪���]]�����He|M����5�����S�/���M*~:Y�#�@�Ζ��(�v��l�t�C�rxi�+��V�n�W �,]"�S��'>�W�=�Xg5a'�\�
ཛD^�a�#�Ӹ\�+�C�]��V�r�y�����n�_���a����L-W�Jp�RbPꤤ��� �BsPę�%W��w�+X0�ZQ��d���\���6����j�.3$�_k.xK�lfCĩ��F���y ��$Q$��Z"p=:�|���o1�.K|
���b�X�g�0��A2����C9���X���Y��U,h�0��-7�W#0D�m�j=dx�eQcn�m�]���#��wO��TXGBGJ;`#��^r{�0�A?��a
	���Yf�`h��X��~ �5@��_��3mb��ո�+�t3���[0�)�D�E$ +�sp҇g��&��,��rk���J2kX�Z��p���t��1$�@q���2�V//���g�>�4�,�ȶ�}��@�8L���G��).f���⪟��9��,C������/�"��!�_�/�p��@ m�e�	�D��ꎖ���.F���ŜEck>ο�.��S�^��$�qp�;Y�ٗ�������u�ႿX��T��ܡ����ݬ�{�?����P�#��ؒXeiERk�f��zFWnr��eI<ȿ!?;�b�����f\��*i����~7]�(��Mq\�Z�arw�N�����s��B�҆�{��zh��jؤ�H���k�@�F�rދ�
�������o�'h>�#R|�M Ԧ]dV;�i���v�[�?4��2�=J��*����>&[+;ߪ]��h���@��4B`�L�O���k9=��o�����c�xˆ�!iIG|�m��T荫���W.G��aUW}�94{A
O��"Ր�d3W�W�F�3�:2�<�^@f��NR����{�iQLxEm����ˎ�L~Pݖ��n{�d��,&�4��A�[a9�ZU'�������:�+�<�8p/�ZL���Z#�(����OM��p�m�dA?��P���Q�rf0> (����÷��S�ƙFZl�,\����v
s:b�-��̼�hK��$B�R�g�]1���n�2������Ԋn�'��}��5��(�2��2�>wϽ j�s ���K�a��Ozܹ�M4��E��<{��ط��:Ғ&�����T�mߑ}��Rk
	���Å���F��?�U�B��2�� X*�~� �ƘY�B]K���K�v�Te������MA�@ݔ"9l�}Bj~���Q�ĺ;����s�n^��5���x��z��-V���8@#�PpV���2��t!�#�X�S�yN�푌mJY���f��ԙ.�D���D�s�Bޖ�ZK�ʜp��k83k�h����x^�P��R76�	̡F�C��;�.�c��{3��N^�f-�Wc��&���dӰ��$/>6m�q����
�{KF�D2��t.��g��C�
�e�Pi�$(8��*��"��uMy\Q󈲅B����4�`�|���#Y/{�t��;�<A\Ô>iz�
I�#5eJ���]-���
u�L��/?eK�*۝j4I>([� e����D����Qz;`�Łސ"DvQ�8:D֫h�s����� {��hl>տ��(4!kJ�=�N�:!�-����Q$������r�BS�� U+*ؙ�ڎ�a�Qih)��l8l�趌��NȗT�<a���]��������4�xDw���}9�9)>�s���-��~u��_����~v��yimz���V|}��`g�f'�e$G��!U�C��>&G)<���:[��o��W_�_/ĺ���|�u@��X��G}�|/�z5�������u�T�ţ-W^�E�`�`�̯�F�"=�lW�0<�E9�f���T�G Q3'2J�*��^C�_�H��� �v�
���n��pTy,R�DEj7(�[Ũ��y�{��\��Y܈rA�`h�Sb.�F���A0��>Ap>��\��;�̺�gj7�6~-�tވ�Q��NEt�������,�d�*]�wB���Iv$waH�S�w��v|`��8��k:�c��@���}��?7C��3��}�p#�P�x�B?�ǘ�ƖL|J����\&�uYŴ�u�pz�����B�5\?�iOo+y�Hze2I8�*��X��ſ�{aկ�pH����,�� H��}�-z
�P�LR$"y%|��4�g1�-M_�����ڤ�;����4=�a'�wgM�MR�&�ب�~��y�����9+_HYM���^9�� Tm�����Y!��^Ui�ϬTt�ָZ;	��{%95�$��T5\ʏ9C>����(=�*�:�	�!��R��\u��?�#4 r���O��6�:t��Cuk���ǹB��zjԅ}C,��D0��A���R�AI��~�B|�P�x�T_g�mJj}�C���`�-
�M�Xl�����;�v�Y����:$3C|�l�!g�nT,�C�@^E��؜m��@��~�dfGJb��z�2�f>ӯ%���	��C&��ixp��rE8%ی�\Kл�'N�b��]�ԍ�QQ�w��TF�ÿ́	V��p^t8��O/��o<�w:��R�!���W���c����?�pϻ�Hb�UJe'���{���ը��v&�ؾ$h(�v��-0gO	YD���\׍δg��6��i���
��q�dV'*�|Ll��U_���;�����H!?� �|�"�����BqP獀%�/�nʴ��q�X \���'�.�t�4����q��\�A-�U]���Ύ�;:�^�sD��h7�V\�R�b5�� {����T������C�EI���Xf�7��X�n�˚0��m�������V���d�w��w	\� 5���I$*�Y��8�=Ir�s����:��<��8a� ������v�!d��0����.�F��n�{�HPנ�P���F�p��<2K��3]�\�Ԝ�R�K��KT������.K���F�v��!��4�]������� �-��"j����Mm|S�߯8A�~q�^?_ۄ����+��Sz�'�t�r󧌊 \̑�U��G��'a���Ѩ���rGj�|�,5��ї{X�X�L^�u�~�a��+�0���r�V���TXk싼n����;��I�tLH��J��b�^5���Z��.�sK)*[T�2wiX'��Z�G�?J�=���e6��S�u3��Mg&_���.S��lRf��D�bF�~-ygZ��s��$�!s"�a:���|5��o�3Kw�Ӛ'�2X��0��2$���������"z�j�t�h�_��aG70�*��dDX����s��Q�IYm��y�B���0���eT�s�G���#���r��o0>��ԏ
����[Y���h��K�
O~{�j@�R;�4�z���ް�f�5t�G(�V�)��E��Ԏ��*r���,�������J��U�~��u�=��m�OS�1_��@��-BV����ۋY�(��2�k�t�{>�L�g=�Bd���!,��ڪ����fg���.��*�"L�v�is�J:)�[/�m�#�	%����}�ɨ�.���;�c���oh/�.̙�$x}W�6������j	ń�?K�:�<�/���O��_Tǫv��{����'3��4E-؈�� ��(�nm�n����za};����?��f��̤����X!�~2�رi�ͼe\�Zb�rR��Zc���׉�������W~h��jSUr����@�Ȧb�Fcm��T�|�Q��_o#S>̎�|���A��V6����`��u4��2�ܽJ}ȳ�����L[&GĪ�42hgw@���B�(}�*M���ؠ?ӿ��C��x���<"�G��i�4�T#u�2sY.B�ao6}x'�Oo
ʴ�"���dnI�W"�:3�������@!����kG�͵=�i��x�~���ɎL�CP��-É�������,a��+Q�V"�9�u�U�X���}��	�q��B�<L�/s�����Z~�U�	�����I��HrAz�P����L3f��?(�s������q�t�$��D\,�qn:�E]-T������Q��-2�#=̠��i݁2m���~�ʢ��}�)pQ(:YV�,�>�K ��%s;����B�g�j��6L45o��5�3=���U��U�xH�Gh��,z���
dH�~ @��iz�JUAU�A�mY �a~�{!S��bkK�ˬ��b=vb�δJ�0Fߊ��s`���C�O��l&�j����l����7����iOY�bEh�X��x��z��-1���s�gس�DVȺm�wm_�/��#�t��Ne^ǌ��<�^f�\̙�-�ٸ�D��@BY#�Z&�䜫����Ck����i"�x:P.��R����E�����|%�.�����i����lEW��&p$d^�yg>1U�q@��k������a2��ti��gJ�C��$�xw�P$Z(S��*rf&ݞ=�y�ǈM���e�=r�`�e��#�/��z����<|*X��ӗu�I��_e/H�x3�0�
��TL/�`? LI%�ij�܌(� ��/:2��a�{Q���`&1&ދvv��p8������Ji�֝���bl٫����f!�3=����U�2ʨ#�f�$��,�S����B�� �iش���		�,3�)ۻ�8@����N#�Gg��YX�=�Z��n��o�D�#������Q)��:\��(���ͫ��5���Z�t?��6����� �Ⴑe��	��tю���&������[�!�m�8���=���S6 �p���kCk���|']
z��ߒd�԰�ǲ�x�(���\���v�6偊�78=�8�>w���g�f��(\����3B6E��!�^_,���A���v��v�J�&żg�ThR@j�X��"�S~={�k��:�V�-ľ`���b����L�|���ٰ3>�w3ַ�ܘlI���g�T6Y��t�����N@���1�#�~|�,�*�c�B�8����!w��5S�pޢy��`G	M8؋(:�������ؘ��ǎ�N��pޖb�{�?-��?�L��i�E�&��[Y #�uH�@�:x+$��\z#�O��5+t4�z���8i��56���GŚ�aZAp�Q������GHX��H�T}����J$].-|�S�/t115M���*�B�#�#�4xG�'f?ZHO�RA��:�:��9���t�9f*H�#�*^��� �D�����,a�9�k�
�oT>�ֳ�[	+�%��b�?؝�ϋ��j_n~���&�#Y*f������1���u��Z�� ��J�;6C��cիkʊ��4d������t�,�f�?��3�չp�\�l��T��?���|����W�3:��W
�{������M�*��)���-�v����+r��V1C�>1��4Pn��;�~�?�dm�ӯ��+��տ;�d��bG��z�Z3��a������$�+᜘@��p�SSr�~7%�_���y�V�SN�T����a�l�wM�Fb�߄D�h�yѴ^o�ȑBC����<��Q:R�Jm��I����nc� 7��&�p��
H}��J�kI���K�.�����&�Ծ���1���H<\O����\�F�D^6p�ia{���
��h�0�*f��l�6_z�;㶦��bH��? 
_s"�X��uKq�W���Q��i5u�N<VX�q��-�Z'���O��4�=\��T��bA��]���������9	Dy�7c���S�b��" 6����8�7�ѭ��I�XY��$�n%�0�����r�����"d�(rd,���r���CI5��h�d�i�&�@I�T���od:w���P�;��og�Q�!�i�0J���)<F��GƮ{�\���]i��@�<ͯ�.U,���ɤ��F]�~ȏ��1����L����I�c�MN��FR���]����4����冕�)���fWS0��T6~��弙.v*,��$+�,�d��t�t�rn6��-1�̕пMX��"���<2�s%���-����5�����oZ��r�^	}���w���+�SgV�Z���W��&��n���s4.���Lc�MJfG�bԍp����V�OsF�6����&�XB^JZG�$ߩxʺ�T"�6���ЂĐ����t_�� ..5�l��g�߱�F��by�Ԋ�.��$ȞS"f#Q:��|p�&og��Kr�����!Xo��0�p�2�<��l��&*+��wu	���իh~;��2�|7�]
�;D�B(���jnnBQEem`�4���m2���eTο�G���#�5�r1�0�k��
�a?�Ǫ Y�&h.��~��@`���O�)cqYދ�l�#�ti�)�Q��)x�E���ԩ�-�}u���P,4]������"J�H`�������f���*0m1�X
@�t:�(�V峣Jܓ�tn��"`i�Fmz���QL:R��=E������[�&y���I����w�?���<I�%�g"�&L�$�Z�e���=�m�}	`W(L���|�.�n��;�hc�J]�����	��Դ�$�v�1w��MfI�%Sm��������
)������9�qmn�m$!��]ϐBp��N$E���-�d�)�nh����5��;�����."f�M���x���~-�����w}\8ZZ�L�r-B���3ݧ3�X�Ÿe�<��p��h'��j�%���h�}�A�F�C�Au��7�%��o�>*>�W|(���ܘ}V1`��Co˥�z04��$2CJJX�̌u�t!�[!sŪ�Xh"��@�
BV���.��'��V���B�p��xA�p�W�ZGr�����T^|I��a�.=G�a�7�}3Tuj�
E�*"���d�[�W���3�4M����@�7|	�=��h͐Yi�4tx{����Qd���(PS��ä�RZ���d��,��2�ƀ�QE�9Y�*U�&����u��zQ<?�/p�Z�;|�b��t�}�o�#U<A��P$�f�G��f���(mWs��M��I0�OB�7�\ǍR�l��H�-�Ѽ����l�k)�w�g|��d,;2����g���
���J}�fb�a�(՟W�F�>-b� �S>sV���A���BMK�/�>4� M���j����,�p����SGK��-�ǖ�����
���9��\V�Ŋ�Ua��� ��~��;|-�ظ�K��z�A��v=T������玼�[�5���
d�l-�Ojt_ׂ����0H,�0W��d`��u=��ux,Ukzu�O-~ɮb@�N�1VÖ���Ƞ��3#(uzI=�N@﬌����8�f� ��յ�
~D�e$B��:Z$Ϝ�O-��U�k�,.����x��|PIPVR-������N��/,.��;�1��$� ���WYb�&K�wdI+���7>,]�q�p�&�h��a<�)2dT�t���g*C���ө�Pߏ�(n�*�>��y%�y�����������V`fn��D�/q�l�]A�<�a�C��p]	IZ
e��C��#��AO
��qLj�%?�l� #Rj�{(�8w �����'�<k�Q��>`��ކ �vk�8�w嫞vi�m��x(b-�0lt���!!=~=b=�p���#s��A1�$8H$���|�B	  ˊ���=�ڄ�:�d)��8����L+N~6��/�+��߸�Q��g�"�D��/�������ɤU��U��H�q�ﴛ�o5�0�����1²\��e�ҖDQh��W���&��;�[�.[�iڷ����j��0o��k8���N��J�|B��z+���?����qa�M�d�#���^�4�։P�Q��<��=�$��y޼�{�=f�1~���~���3]Z�� ɪ^��蜾`��6��v��k��g��w�T7wrR�	Kjʚ�џ3��|{�#ʕ���f�`���b$�d��ٱ� �t@�>�� ��z�'wIeMg`(�64=�tT��̇ӸN;�L�� ��95�,4�*S7iB]{ʄ���w���S��0���&`M�8�F�:���މ����u�P�r�$Zp�e�!�?�z5w��L򒎤�J�&�R~Y{�u�9��߫�7b\��"OHBT+o��z�.8$ԈP����u��aK$�p~���1o�HȏH}�c('�W��_S$�I|AУ�*��1r]MՃ��E�ښ���h�4�'�''C*�Rj{�N���wq��pd29�vH����a^�+� �U� ��OX.�k��Ey5T��֮x	q�P%�L_�Z�-�Ju�E�O�����9R���*�A��%�!/���8us�%�� ����E��6��/���k�sLǯҖo������,e��:�G�wD���r�wѶ���������t׊��� p���o��p��#/�M~0�d�*���iv�	,U��а�SC�蝟"Rn�m{���r�����u��E�z�d�Q�b�0#z��üܤ��[I���چ�s��qp��r;#%�RX���Y���wN����Ǐ�JU�"w�ZF=����^�Rv^j@���V׭lM�<��:�(RRv�є��}�4vc�_��d�pE�5H��%J[�]����H���"Oy&�,����!��ch�O�����u\Mb���Z6ei�v�f*/��Z+�*A�Rl �*_1T;�vъl[�H�t %a�"�1���j�q���[�
�d��&dX��b�H��'/�*(4#��.Wg���A�]hH��:^��1љQDNR7�k�t�b�8 �����������|�IL?�X�1���n��0H~G�5P�z�έ�!��d�ޚ�mcp�Q5r?��6������M����a���:r8R�R�"�V������,�~!�;L0忸�$hZF_��>�{*�ז	�8���<h49�)m��H���V�̠��e���~�����祔�� Oм�i���ߪ*�J]g�v�ouB6,v��^�F����~�S'`;�.��~˖T��q�Ζ�&ɇd���t!5�r�늼{���߿舨�ɰ����.T��3<�rT<5������^�Q�4f�����+,�3��{�Vf����v���0n�����M���*GL~�J��b�ܛ�U����sAS��6Ď����X]%JZ�|�������l6����+�_�Y9Xk_v��.	�bl��G�z�zF��Syo���u$�;�"�c:�9�|��oymKm���RpX*Z0��2Ȃ�G԰�a�X���s�*�+h97�M'�7&4����DΣc�;wi
�Qt`m�4�Oޫ��S��*T	,UG��#���r�9V0���F�
z�ƽ��uY�!h�i:�N~1zu@l��j�@�(W�fM!ܥ�t���Lǔ)ӹEUQ��
Y���G�,o�B<Au�܋JC�F�v૦���'8�-1��N@B�#H�V@�����ch��k�!���d\L�\#�8�:���+�AY��-���(����d�j� "�"o����X�����Ql�mp��	�<�,���p�.W�����c� �e;�����y$��ͦ,6٨���ل�a��0FL��e�R�uϕ��l�����s��R{�]���3�E㵔�h�"�KKZnc`-v���@;�g��5�f��ݤ5z��(~(��&�2�\S��ZX�@r����#F�Φ߃���җ$%�+cShB"�jI�^菹>����F��ޜ����].1�oz�>�ā|c D�wf�V,�D�����&o4� 92���J3Tv�V��Z�[��n�h�Ğ@/��Bѫb��.��.*�u�T��}���vx�k��r�OG�E]l�T��V�hpe.8)�a%Y}����
�c�"f5�d��WXS33�ᔂM@�c$\�a�d�k!�ir&x���~ɚ�S.P_rÿI�դ��?HM,���aйL�m9���UX^�)���XD���	<zҽ/�*M��Z4	Y��� ����Oѥ�W�A�z�P���B�lfA�?(([������#�*�i�1\b��g�Kl�-�J��:r�GAC�����x��_�02#)�"���%�ʘ�}�jk���(p���[>�� J�:sq
oϼ{G���j+%4k������e�DFs������m�.�^�r��b���b
���U��2nڢ@�U<���; )��~��'#�s�K֥���v���2\|���3��l��4�lHֲj�J�����k�����	�_�;�ƒ��4uxG(Vz�ܔ-���#���6V����-D���uD#C3�ľ�N�B�O 䔌df��o�?1>�O|�DPBO��Z���!'3�<mk����x���Pd�:R���	��08��X#.�ƌ�U�߅���JnW��.&&h�d�����>'�*q�2P��M�Y��@�2?��t߄0g�)C�Ғ.�P�-�(�:�*h7��T-�y�j��e���%��L`!���4��/�-K�8��<�&ޔ�^�k�I��4e{v���N�&Њ
�.L��~?6�)wVjEc
(�w� ��)0�۵t)Q+O`\hށ�vbi�8kA���w����S܍h�l�o�!|f�=Y�̋��ʞ���k$s?W�6�1�Bdr� �j������]���&�)Q&68=�߶}�hNٵ��̓F�E�3���v�j��rKDH)��
���J�'���p������m4�H�;�O^��jK���[؇�]�'�K�י>e�����&�Վ�`&X�����[�웷c��� �k���GO�f��!z��x�)|]Kz��7�_p�&���軈�\���g����lw���G=�0�ٴe��%f�s;��>��x��3x�s����^Ԭ������ѫ�v��ܩ L�2��TR�aR6 j��]�=����S{��������)�`���b�Z�s�����d���>����m�X����j�g��Y6�xt�B!�"�N6^{��-���9,O�?*�*�B8ރ��Pyw2yxS��~�/<`��I8"�:�x�]
O�8y'����v����pTTr���?#�R�kL-gg�{��&�!�Y�_Vu�}T>.n�ӛ�\��=O��+jH#zv^q8��&kN<��?�P�a��p�C���J����H�K�~��s®�l$��x|�l��%��1�A�M��D�`y��Q��u��4�'�'�.h>%eR���	:S�����	�Kt9� 'H*E����^J� P��;YE�ʣ��%����oTEٛ֩��	�k{%j�uƲŘ� ��\�\����;*��:l�<M���uN��:H� CX}�@�6��-��Xek }��*@��JN��6ì,���5����u��KSY���h�}#����3a�%�\��C�{̴�tؘ�O����MY.����c��v|�0�}�k�CͲ���/ n�*��+�/Z��5���o�5fd�b=�Xz�
�����U�����{�����p.t2r���%le$�6�Ќ �N����nϏ�i��Ew
�FS���a�ܯ�O^e�Ǒ����'�<�yf:b�RQ��52�ρ�c��!�P�Bp �$H�R�J�T����]��,���~&)�5�@�����~�~OzgL�_�\���8��6	zi�h�!jx�j�EK*Z�l[I3_�}q;�V���:�HR? @�{"��eթ�q������_k*�1�XQ�q�c��'��S��4^�ی�y��^A>>]#)Q�UV[��OﻃD��t7���ݵ�bFz� �n�ԝ�-\�Ԓ�I��X7*"ֻ�n�O0u��P����Έ��<�	dbB|�h:~m�5-�cĚ���h�ɹ�����N��:������q:T�e4U���!.�0�����F�����}{E�����͌�!�<��$�"�RL?�͜�l�t#y������O炵����\�	�w�ɨ�4���L]B������Ѧކ�,=��~�9SB�E����~�Y3�:(��i��6����X��t<purd#�����BȂ��ٰ�-������R��Y��=�5�#�H�z�)ʶ^����t��H�s+G��I��VA�Q���\��n��ء)���z��L��=J\&xb�K���h���<s<�(,�c�:Xx�Z=G��7��Ti���x6{"Ά���^	T*
_�F.��l'\�aF�/yx)���{x$��l"\ĕ:���|�o�K�Kh�}�88X��05��2�s5�"︁��͐��q��5���+h�R �h��7�*����D	%3���dƏQϛ]m�8�j\��c�	��vTD��G��#�# r��0oH����
�Z��}ºYR5
hd�5抠|~�K@�(&��L�Y ��A�Ht����G��).vE_���I�s1꒹?,���ו���s�J�������+�\���I�1��@�ӡ��eV��_�wЋ�x���:���u�,(�Lp�Z�3!%�P�R�_�\Y5��0j¥������G��k"]�v��n۸����̺pmK]	���^-ږ���.�u��c�֌�����y��J]7$I`]�'��ú��F
��"8��*ƚ���܍���0x'�g��#צ�<g�x���Dc�E�Ԃᣏ���Kn^�F��[ȫ�P;�A��yf��~�p��)�"~#X��zeu��7\n>%ZӷVr�h�4�i������򎈐�$h]��j�&�9�y2��w��F
����p��*�I�o�՜>]�|�&8�TwV'�ۉ�� �G�14DU2p�Jʯ���"��N[+�ɖ�h��@J�BL���O��Wj����+��&��x�M���Gh�%88�T��7��o.3+�a��W}�B��h
;�"A��d�W���3{�X���S@RN?KI�^��FCMi=��x��k�yam�]�SP��J��#|P����,d��?hG��9]�U"�DmH�z���{J<�E�/DS�ЪZ���t��;P;�s��z�A+�ZPZ'��=�f���(�~u�/d��?>���X*\���bZ9��9-��f���$�FҾ<RS���X�Z*b2~~������@���#}t�D!��(�b�	�=>�t3 �s�fh�7[l����ܥ��4�4��K�D*������^v��˪	���'?��/���R
u��ȯ0�M���UTU���- Ĉ�~�L�2B��.43K��n�7D>v������*������d�݀%�lc��jjVC�\}�Ħ�q�fr��Z��s6h����xbIzk3�-©��$�؄�SV��S���`|�#^�?`�N�p��Y; �/ bf����f�
=D(��Bʈ�Z���\���k�p;�z��xk�P��R#T�u�S�23ǰM��.��p��佈�-����NWOG#&:qd�%"�P7�>"�AqQzP���V��2�2.�t��gPI�Cz�C��n�PU�(��**�O��/UyH;�������N�9`����O��/g��Ǭ<-UϔyT�f��I��e6J��ə��~�
��\L��k?���vj�V9(G�� ��������Qf^`�3d�|^tv��:8&+�Ԙ��i�.���aIl��'!ׯ�=�ͻ̦��r����$��ZZ؂��B��Z AjA���z8D��P�)���8���xlBN4U�x���a�8߮�C�Q��� ��D�p�i������
���cТ��f�r�p��G��@��e���:�B?�B���RU�e���=��K�|aU&��;���2[��e�ޱ�|��Ħq�$ �a���|�_�3�O|x�'z!B���ߨ�a�>ǃ���w�_[�L�P���2�@=k\+���豳4f��T�9�)�3��3���x~^��2�4��l��v��ɩ[�����Tm��R�N�j�~�G��$L�{��#�Kw��^ `��;b�3N䃱-������>�`0���v��2�8��gV��6��Ft��̽('N1셁B{��,j��*I>Ba��5/�w�S�ɢ���`x4�8)�:
n��88O�sb-�������_KMpcp���Q?���-j�Lh[��"�&�xY1.Ouy,o�騟��\+�,O~�+e�z�W�8����
��+�sa��p�9�������H�����Vd�L��w�$�|w)�� 81(�MKٶ�{wڐ&��PRa4)H'7V�9@�R Pr��E��Q@�;ĝ&� 9L,H�ך�|^�V� �M�V���E��� ���T��֤^�	'<&%%�䴐qf�@O�����/\����.�m*wV��Ң�W�7�	��u)��u�@ �+8�;S�6T���J�k��ǥ���%*��qx,Qµ�0���-ǳ��#��ق���g��s��<�A��EI�� i�Hr�/E��N!���M4`4�ډ���͍vw9��2�&�C�o�]Zn���/�uʃd�Ĩn�<���4)d��4b�Zzi�ԼR�௑�Ƌ���<yA�qL�pI4~r1i�%G�`�H�j�'V�N��<��������=qw}�F�0x����J�A^`��S�����<�-:��XR,���p�t�j��c�}q��A�p�"�H��JQ�j�a,����{�X\�&��M^�b��� �O�V'f>�\öh���6�pir�[����4dP�o*��l�P_K�&;�V��":KH*< [��"y�Մ��q<hT��x��Z6�_[@Xs��~�H'u�[��Ƕ4�o�d����2A��f]�)0�pn�'���FiD��74MZ��b��� g�����j�����I��X�BKֶH=n6� 0����k������ce�w��d�ŕ�c1��f�5�bĵ����{ڤE'���%n���U�:(���+uЌ�T��{n�� !P@j0S��bF��x�k{`E�׌���\8�<��:�������i��o�� �x*�75���.����3=�2Vm�1vR� �]�L���lA�������9AS] 8�$O3~�<��JxSG������=�$���tW��r��z�rw�}��Jћ���M���2�ޟ��hG�5`=Zу��ĥ�^�	�����+b5����V���@����n��M���ֽ5�L���J�ŏbe�¤�җ�'5gs7�D��ɀ��X��Z�1��q9�)�^�%6v�I��0�����oQ_l�k.���l>��İ�sF��jy���_�,$֥"�D�:`9m|!�o8>%Kc(Ě�=.X��0Pi�2?���)1�׌M��0������h���ۃmM7A�jmDDƖ�q�_�`Q*�Im�����d����c,�Td�GQ��#��~rB&=0*�k9
p��X��Y���h����D~� @�����������ZR
Dt:���B!o)�R(E��)���G��s��mK�,�d2r
T��{�J��@�����v��"�����1K�t@x��ΩV��{�T�ŭ�瓉ն��k�gnL�i�.�����wyΪT'.LS�K������L"�_��U⸶�\�G)km&[�	�G�M)����.)��l��c��`�[�q��b�̅a$��$�"<�^���V����&/���mL���S��n��bk��~๸����t�����E�a�ީz���nYj�,��f��;'�h�+�vfel/�����ē�~�����ͨ��\��2ZN�r��f�Fd��������M,���8hx�j?W.Hι�m��-AF{��R5:�h��d!oQ8>8z'|�l�ԭa�V"Cn�T���x4�y2~68J�_y��E+�[�q�$��hS��@e6xBǮ����㑒�L���������3�xrO��FG�>R$TR���..M�a���}d�~��6
���"C�dZR�W��3v����@=ZZWQ �!��ixL�xL��t܎���P��G��������,M춄���Bn"9j?EU�O��_RS��IG�V�j<��@/��0�HZ�1�,��V {���X���HAf�WP��/�8תf�@(�¼�J*��+e�����n\����]>qn-@�'�g��=�uҙ�n�4�8���U��2���S;�[ �ʎ�]}O��\?�(�3l�T|>>.A ���s���ϲZ��ӹ�����4��ܶ�U��u���ų��)��䴵�3��ߘ�z��b�
�Ř�j+;�h�ڢ6�U�Z��Y܇ _ph~�' �|?�鹨K ���$,v�Õ�6���i��Kv�F��;6�l~1j�ۂ7����·0�US��ƽ�DL x}.Dz�C-���_C�ۈV��-��%��R#y|�!�N�a~��G��ʓ�f����O�ſBDC�BE�Z��n��5��r��k�B̺է9x&N�P�l<R��CP(��mUJ��z.�4E�B!&�U�c��W��&�+d�RU��:>5�q��p�W:������2��EtU�xg�hCu�p�� oP��(�D,*^�.�
��y�a_���0���30�y(�2��so���N����@��c�{��~-��I�)��mQivސ�#�f=\�$G�Ѣ���Y���}atlf�&��;]���{��R��k�*G�<�g���@e�fp��K�ox允��(��a�
-���8"p,Ś����	���S4>��50��O/RZn߱
C��z��Z=NR�E_�!�^5�g.�s�����1�:�,� �Ĉt�lw�7ZmgCDl�}��|Zu�y~�A�s<_O�tX�hjZw	�(�c�����/��AC}�������f����Q�(W0F�S�7��Y&�B����$(�ݕ���Y�FĠ Em���,���Ķ�6F�)(&�M�������T�O�c"N��<��]��5H�����v0P��G�O�h�B�|����3ԣ�ܕD��34~��1p�i�n! �`jPC��j	_��O���N�"nz�HM.��63�D�|!�(ȼ�@*N{����o����8��ݪ�6�}��AH�9g~䐧tJ1|f������'�˅㔬�]z�➨�@��狵�?"=W�GP�r�(˲ME]%{"�<b/��o.���7��l��{�Zp�O��������DB�e���7ƌ�<������n��-�_ �#*D�Q����[���<���5����~� VC�8�	8b��s���t6�j�0���9�M�5�i�i�ހu���-�̤pm�%=w/�����şq/{&����DC���q��'RU�3�R��2 X���T�����g��b�� ���R֓��kdvG����)�|R�/ɽ�&Lo�V�0��sy<��:�߬�!�Qg��>���-�Z�g}�yC���_sK�|��X��S�[�T:.��lC�a]��/�7�w`��-5P�S��_ػ�Q��&UdM�o-5�?n��;`�/ۅ}9��E/QD֍�	��#��-��#�я�2/P����TO������o��d��?�k�d-\5�6�	�\-��Y*�d�ۊl�Ԣ��]��H���Y�n�_����nVFϥu�x�s&�-���2u���V/мw�nA��Sr5�
��!�ȝyIi9
����@z5,�EC#�:�a�ov�ȃ�^���.ZY�Ź��"}�}?8���kZS��g�ufͯ�o��R�E#�"����4�b��=��|3[F��oRf�t����mhF �J�IG
h�|��!@p6����G��@N�7>seIR?���!�v&�k#p�$W�M�TQ7����ɦ�0%�_ѭ�\#�4!��!@u}
4�������>�#C0��U\-�B:�!W��`]�kTf������]��q���Y�׆��XD/���n���8��;0�r.^�Y,��܉E<)!�h��d�tq�r����/�T�	vAvU�	>ܓ�Fl<�3l���O���k������z[�7�>؏e#��P�
�os3����9�(����GM�݄�����e��֦$H����.�(��*�&����S�ţ��$e�r�*�(R79j]6ƅ�?�dg��Z\�#(W��p��G��N�L"G�mN�+?5	�D����DO��<Y�P�7YpLL����=~�R����Ɨ� ����^��n�&�jj���2��3���+*�Ch�q.׍gr �����M���2xUX�E`�8ω����'�l "�(%e�0�e4�}��Zwk�;E7�������˟p�����y��(�EEZ�n���?lу�e���AE��ZJ��W��1�מ8=N��<�B���S2 Y���F�9�%�Hc��o��5��\ƁOSf/�F��[\̧\ʴ�/���| ���?��h[l�	�T�[%a.����cl��75��v�w|h��6�{��AY�K�ª� }5��L�����f�?�ߏj���'F���f��s���ș=�?�رn�I=a۫�����霗���H�b��1���e?���vNu���{��sh.�2o�u�:���5���* v�P[T�h�;*J�FТ.�q�_��҉H�gKԯ���H[�{������-�bH4����=*N���5���k>b�Bo/�Rn�`!w,�#��ٞ*v���>pN<l���Y@���q
��awQ��|��X�N?���Q�ld�Z���(q)��'C(�o|�ީ0L?Ȣ�Q�rZ�-�#E���O��+#�,G���Ep ������}08Zf�ك��+�ð �6}���Qo	S'�%C���V�+ڜ4X{^�wLРr�A�}���Jdq��B�Ϥ!>m�gخ���T����r�2����,����.��km�EZ2�X�?C��>T�Gt�U�����Z_4�ӫ;�T���u!U�Gip�L��C��S��S��!
,/�0
Tf���3�^C�Q�$�Ť�^��!9]�f`ay�ȳkrMX�6Q.��� �1�F�j���xߖ��0�Q�:��澀��MN2�~P��z����2Ԁ�-X�<��)��R5]b��C| #���������	æe��U��0��b�5�|��tqK�"�9S�]�¯2�D��|�^42@���GK�J�����aX|�N�-�-0��q&CwvQ��^���2@�[�l�Y��c�Ϡd�&��uS�j��(&�GQ؋p��F|�c!|��P]���-�tf�v=pN$~Zy�p���4��#>1a����P���_�*JvY���,C)��ђ���s�[�NX�H�Z׽�p��{���b`s9���ޠ���(�C��h�F�Zݵ����@�31�`xpEL��.�z�a��đ1�[~�ݓ]j�F���g�+�u���/�ߋ�˝
c͓�cE��@�F��m+� Xm��w~Y?��� A���$*�g�j���rm�r���,��:�ŝ��2�*�^Ub�k'���q�m�"*2��f?�x>�clGf�����c��_���a�5�T&��u��CG[H�Lǰ���k��_!��.�b�T�L���Do� Ń�T�7��W�!+��f���:�nr�Ƶ�(�D�*�殣+��i�
�o��|� <����4À�#"M��,01;�l}w�oF��-
���IF��S�b_�C.���pi�Ϗ��O����G��0 ��b?9o�.�Ntc��8���uX��ĺ�$�>���м�@6+��9��JM��da
�N�é-bX� 0w(z8�P6s�d]�[Z0���c�7�d��7���Fq(0`G��p'3�?�c�����;�t�=b1e~��p5����FJ.aam�ª��_�=����X�j ܝ��혞ϥʊ:�/����(,{��I$5aPE��d^�,$��ig����������$��ɞ���Ӱu����~���߰�+��%�6�?��Z�B�����C~�'O~:�]c����r����:؞�cy\��IwP��X'�7�p����.3�d�ؔo��2�j����!2��?xp�:��j�;w;�v0�ZX\ ���2FI��tD^��㌗�d�n���L���HѦ���7xY[Ur	�ΝW1��Ceo��n0�d`G�RuY�K�YY�+�X�t��3E�54���g�m����.!HӼ@�b-�0�3f�O�/�9���2D9���pN!&{@dae��o�7o31�*�٣�{�{/�pJ�����t޴���sh�p��q���g�LKߠn��e�=� $�@�9���xgQ��2K����U�!��K�f��e�`N��4�H��`�|J��X�џ�.�<��"�N���3�%D`��RT��fIu�.�7#: .�v�M��q1�u�j��è��b�j�:��͙~&�����u%�:���G�eF�^�O-^rй���g�M�*L��AG\�}a{�O�^T����=�x�Wr	)���V��\MtT�Z�����;�������)F��n�s�7;�z�v-�p�k���"P�~�Lȭ���̼��|��)n<y����V�U�P�6�ݗ1vo]S�65��	��ձ�j�aK�ŋ���/�!f&��P��M;Y�>�V8��8jv�(&/|����Ēz���)#��ڳ��'	16�H��;���Rq*Ĵ�iPC�V��K5J<�.�2ed����3�c���� �kQBula�%���~�0�z�O���x�i?N5k*� �z��4[|2��E����H7�xr�}���(
�ai�l��C&q��K�E�6�
�m��OBF��ߠ�>�ғ��7:�䓢ǃv�1,�AM�Km8B$���q��z���B��Qt���,�����
D���<�Ͱ�����`�W>�jL�F�J��ӊ�#��㦆�ӮkO����\}�Ğ��lM��Y�K�X��%P���(�RO����A�r�ʫ����:G��=׭MV�r}-0D�~��������,:<�i)L�|���Ȕ�'����j��挺P��g���/9a'O5"����&9I^�&�M��۳��xO�a�i��e�K3vL����0;4�<�m��~���_� ���ܢzH�$���R;�(��������7L��X% V=--HL�m-)��6u�9x�o��%D��9�;�#ڠ3��Φ�ze��;�pS�Ȣڻ2����@�S/���6��i��/~�0Z9A��*�yp�����`����">������m��V��:��n��;�v�F���/�M�~��&_V�zo;�)WhC���ɰ"2�Q[Ӌ�޵1(��`���@��}ͤ��_��p~�Չ��B 	����
�QT�A��}���B�1�Oo��N�OW�-�QG�
���oj�����$(d���ߥhW�ب\S��^��<1���:Cd�3�	��������x���1Qv�vz��%s8�+���W(��;�ݣйx�@V��6�5L�?5�PTm�T;]B���(�m�&�P�=V=ժyC	�r�GS�2�e��%ӷ6"��s=��%�@��r� �\-���#`r�̟�y�{վ����m�\�o�P*4���Z�2�I��q��,^�׆="��&���,���:�ެ�vk�n��s�0�t���&	�1U�8�!�W�+����!��*s1���b����u�<��M K��}����ҥ��!C=q��ڴ!#�2��M�ұ��n,;��'ׇ���ߗڌJ�?+����D��2��4��1U��r'� �,4�y ��*�����?�=4Q �z=�1I��M� .��O̨$FO�ӓ/�Rt���9��W�2�l�s�.��BȿehF�X��Xc%ۂE�`�R�-i�.��V��[@�f2T�^�?�z|-'�q��B��#���P��zj��L��,����.��jsB�?����T����t���N(������j���j �%2i:�L*jC���'�A�}�.#`|�8~�}Wm{�i1`.�a��;�U���C'�D^fr�?���A.8�'`��P�>��o5CD���=�$�T�i�v^I>WP�~ju[���%�AH8��gq�㵦n��4t��,!S�0-����x����3".��꼉�	['��N��%�X��.��*I�Y2�{_��'u5�w��Φ��y��^_u}�^g���5#��C�~���"}�w�\�?��l8^�~qC�p�P���7��WW2Y1���u�d0.���O`��r؅��ƛAc�-������J?�,�ҳ�.��B�c�Y�27�s?\;Z�op��ǆʉ6�/�d���#�{Iu$�D�E8m��?Cc.i����U�̲F�T$6����q�?w����~��Iߏ��V6F�&�h\�B���
���F�~9�cl�!�TW �L���y�&��CusP�z�&���O�d��b��=������ej-���@�2��zݥ�y�j14w�}vo.��"� �һ2E�a���D��+������7�F$T�
�ѥs�Ƽ<Y�{�Q�M�w1�m���������G�F�Y�������+h��ӧW3��"4�5��j6�L��A�E�iy@�|��3��#�Ne���5!D��\#KN��@���eN���vDM1��k��Ķ{μ��ͺқ��q;o�~���f2h
���p�����u����K~���z��'��_���_��9��xF>�P-��K4���4C�v,����e���N�h����(�o�H��u(0��m�#�\�N�S�3�"@`��
�Ԩ\�*I�Q��vB M�z�Lߚ�P�lu�mֶ�~��"�g�z�Y:0�U���{������u��:v�hG��IF(��Ol�������g���د5�@a\��g}��aO��T�Ρ<oe�6+�)N����$\�t�[k:��M�Zt���%��@�)Ѩn�N���J�z�u��[��1���t�]s�l��k��$�:��\��d���X2U��C�;,�V�i���5���Y#]�bwj��9K:݁����ʯ0�⮬��}#�8��jj��
�|]q$sq(���,孷���<�N	0)�H�#c����R�]�3J?i�� V��5i�˰e'$�Z��֯�\c%��8�:k�dl�V������/0���OV��x[���gkiW���3��|6wE|4��J�x���#Z�
�Ăi�7Q�BUN�Z!E�!x
{�t8����c�۩�Ÿ�ҒH�7���R�΃; ,��M	��L9�$ӿ}q����g�����|��� ,U]�sS �I�Н��c�����(��@>":P�ŤJ�H��t ��j7��>Pk.wP�W�%���K�?��A|�ӊ{eX�I%O�|�+���c�)�������-�r����ۻ:F���ŭ�r��i�4k~�G����N:~TR�HA�L���'|�`'1�Up^�%�W�ٓN�f5���Ca汐"�K��R5�9�<C&�p���Ѯ�O��SaU���w3�i:�}�;sC�<���}]��>j� u�8{��HQ��E��;q/�����L�L��YugV�t^H��Xm��a�u�b9��)��>��|��"�?�l�����@�Q!7pr�#��-�FB��.QS����/�]��n�A�O�sA�ǰ�X�?ɣ�����	�ʡLI�<�cm4�LV�a����i��F�W�v���{%�����V���;�(�hg�������PQ�)p�ؠ(�8���y����}��M�����;���B_����
��f� �@}W�BJ��O�1�ND�W#��p?
�tLoIf��U���Fdo���>�5W(h\6�_�]7�x�{1�����d1��	a^��k���J��bx��1�Zv���DL���J�v��O��k��R����f�_���]��%�P8�s�:]A�X�0��qq�&����G=� ����	4�r��S�L��$`A���e�� ��޿d�u@ߕ3r�����A���1#�K���;�ڒ¿Qe@ČlE�$�P	�S�nКZ$;����q�L�^��=A��&�P�·��z��K*Ck#�n����s8���g�t���"�6H�T���M��m���ef�3*6D�7W�M6���?f+���c�AW�3�Jʔ���L@�m,��?Ӎ*D>�t�bs���3�]�ڕp�Lj�M���a��rt�)'��W��^=yk�DǠjH�/�3���Ŧ�ː�!��������z� ��j��/��q�dx���E~g��+�͈ǒ�� @=�%CB����ۥ|Z���;#��ͣ2'� �������4���(�ӓZ��9��Ckloݙ�_K�_~��8�E�l&����6�8�ぽS7BP(*�q��Y�4�Fr�%!���]�o�j�L2���؄S4��$V[�@�\(��M�3��_� ��Y?v��hy_�	��G[Óh�1is�ɵ�leC�5N�1v��th�@���:�<�ZYBP/��~�ô�5Q�	�z�:6AV]<�9��=8��e'$O�Z�soi�um=��$v�;Ja��������:#�z�N�MW�h9�c�,�?q4vl����	�鱼.򯵻��1:q;������.'v �r[2e���1�pA*���Hq��cÄyH ���ԍ������;n�..a�Qb�/���*l�Խ��n�bE:�oM��na��wʹ���O#*�Ƹ���<
��۷� ����M�w�x�|���l�	l8�Q(l�NńЇ�)�����%���W���+?�$�Q�0"�t�`#c�:�-�+�3,���clS��U��8��g8xA!�a�Q+��~d�}� <&Ey)xF,r�8�.�]�ez��>�)_���sT���S�0���f��������`*-蒏I���:�\C��S�]u��};�ش�����1Pr!p��Ź��Mz��'�:�(9�~���]��F�����Zӹ�-j�fD����v
Z�˓�����`F2�+�;X�8|w�%y��tAv���W��M!��Kq��.o�m>{|��?�ݴ�Ŕ��2��R�,���Dҷm���2*.�?�T>�'MG=E���I����-_]��e�^�li�T=�(u��HG2r�L~���;�|4/!S��♑qT�;������X�:Ѯ�5��L�!�T�f�Ao�Q�r��G������R�:u֓�y��a�����7y����h���TMW���4���?!EF]`:-�~���;�Ub���C���fIΚDӏ�3bP�}үE�0�E	b�w]ǥ�t��dox��
Q��z��P��t͟g�_@��ɉ�_�J���&��aeN�>�-�z�^w��8��DwΛ6X[q0%�Ac��9d�)u��E����(o��G�'�p>E��I�c����99��҆Mt�5t=��~�!�pLъ��W��yNaҋ��Y,۫uI=D�Ͽr��ӵ"p�O�U�J�!c�/^$��ֽ{�z�$L��E�5���t�i�6S�M�/�=����C$���ɕܞ���@�g�~�2��'�1�<��6���� EDB�Bˢp��`z~���c�(��Q��c�صkyS:�����PX�^�����f�u���u�ث���)��j�e����2-t9�Vp����jɓswR3�vr�1ٌ D\02�[g��4KD��w��6�{5(��A7��J�����=H�^$�Y[������Je1�<���%Z�� �G ƽYB�����+ �k3�3�S4���Do������w�G�@�]��'n�3=�U��N�R3D�i��VNX�7@{�_e�OH�s1O���p�{f�O�+�3��	��ޫQ��b�.h��������Z�aK��S\�������<9Qw�x�5������qQ�l%��0�=X�eT4�N�Q�������!y�o~c� I�`C����N(��35J0`7���rl����Il����� �H@�����vu9�(�JE����):�A/�5O�$\�=�u|e:r�G1ڍF���O�s�pp���kg'�p
��4�\*��}X�O���T�G@��c�βq)�2~��L\d�����3��M	��2	a�7)�c_nE4D�N�z�!#_z]"#�{���*}�����t�K۱  MP��Sb�U �z�K��~�j��5��L��q����jG<�K"����X���mA�D���Z8�)�j��dϟ	�|�c��!ĩ�.����z���� 	ȭH/;�S��R����Z�iG@V�`5G�cM��Vۑ�q�G^�c�M0��կk(��l؟?R�&��0BnO��x�"�E��kR�1;����|��
Eq3��x�w���z
���iR�C��9��҆E'��
n�V�9k�ҡ�]���*E�7�G���^���,�L*M�<|�G/$k�q+���n��0u��2x�,��t���S��*���X�a�{��k$>�?��]]�J}�9�a�K�~|ʆr�Ek�N��M~�H���P��_Z�"��X�s%�	Y�1𭩧������8)?r�v�ш�:��h�폭��r='�G5~��{��,�|�:�ğ�`YLP�K��5��?ȵ�؇���q���@�a~ܭ"-�q��e�9@��&���nW}�ik�O�5�a�]���xJ3��_����;<U���2���� 3�iDH�����D�;�W��>�ݍr9YL*<���Vt:H lm$`���69/�}�Q�h����ׇ��.���q���7p
���qJ9��Z�%�SB����8��������縧AB�d��Xz�;�������K7�����m̮�V��@�"�^ɒf�!�,�&g0�$r���V)��;W �h�Q��MYz�9��QR-��Nj(m���m�����}$Ѡ��Rð�YՀ
uB��ܡEt�
5#���}�4�B�/O�RGN�w�W��l��
=!$oᥠk�{�4jbdׅ��IW�&�\�[t�����O�1iW;�q��d�F�	�|o�uB%՚eC�0?�+�V1�>Rv�p�<���")��sRFľ��x�GځЗI���Pb1���6��'W����]���k��	�&)�g��=MȻ�P��	���r�֠Sy��
p�\�i�M�g�j�׿��@w��rxl׉� iM#�ap̶�R�rn���+�$��y�P�pw��;Z�h��`�q}@I^�v7=��&<�������-m���o�k��sꎾ[s���tx��&�n1��W8�W𾀘s!���s���5Ŵ������M_ }�+�)��%���9C�pq��K�߻��M�9.G����n�J�'��<�Uu��#��?�آ�EċiP�4փU[�'�B�,��y�q��]	8�v�z4h���q����qq���u�<7#EJF�F�Ӫ=�Rk�w��F��*�S�sx̠�E����o�C�O;��Y�`��- �;�kR)�$�)�'�7��Q�e��槸�3�]�ߠ��OBO�]�:T����M�u+l�����Od�1���̀ "9i���*�T���a�A�� .
���T��r�W�%ti�[$��+�;�s��~bC�}�D%����U���o�@��'�KP����C+&ȖHO�ˁ�T��Dj��^�TJP�]�ubq���A��2�`�j%y�I��{���S7�7�)�p�>xr�#����3�[��x�[nk�u�c%�J��!��נ�I3�7���юÿ�K���R���
��k��uDj/^��WV�m�L+�ݣ�<b"���C�묛�h^*u�Cyw�p����͸~ICY8ִ�\{0������[�<�I��Z��a��T����J&ᳩUڥFK7��)�b�vJ��CW۫V���_r� ��;֭�w��Q$f�PÐ`�l���T�_���d�x��T�Rli9�m�Ul.yg��N�<���B���٬�'��J9���~n)X.��1o��+�����q���
M�*����ݺ ����LS��3c���e�O�$E��$�.� dR�E�������jjz�э[�gP�_ڈ�`����󾐤���\H?V�zA�`�s�k�K�+#ͼ�×,� ���X��tp
j�X'i��/dbЃ���tny�p5f~��E�1U.�я���hج�B@sظ�L�[{&ئ|�9�.��*ɒ@��_6�j�=�)�3�{%� $�͝�p����U�pԖ��j���W�A��=y2ig⼵*�;ʉU͈�{��':~&吶/��^�M�A�J�G�����h'�%Q�<��]]{/"^4k%�-���C̓	���ʺwO<-�i����/JF��d�����	���NR�����ZY���#|�����S{*S��������DrƑ��㐇kh���5�5��
f�����y����ܴ4�H��)��w�J ��+�/��PV���J���`V����{JhlϯtV�\fK&���e��E��	]��[u���}<�`^�(��Sq��2���lpIldv6Q	�������_>q�q#���q�C�ʦ����K��LՆ���ؐ�H�S��/��X����)�iK��������	�\��6%��f���X2j�}������I�5����L1]%��.��m�XT��ݳ��U���m��#���}�ěW�cz15+-&2�����Q����[4�� ���u^�X�p#f���}��}fg��6l��(j~GD����*� y�B?o�{�_f�{K{I�x@�T��[^����a�i��  8]�`v��l���+1�_��j�<��R5h�ECk7ҩ��u썵��Rj�t_��^�*g	���7OyF5 ,A-��̩�t�	[����gh�l�����t�?AO9��ts:�����Ȼ�ʹ��b�/���A�m��i~��qߒ�C,O������:�����������]/(�;��B!��o�[�Zm+}~,�����6�@(A5�Mi:��8,@Ă�k"cFx�‬�D�4�7i�Ɩd]Ϫ�P�/�꣝�=~J�Vl`3���ܰc3��6�ϧ��ԤU#!�0T`eP�LK)j�[�j���K�nU��Mi*|6Νחw�ө��u��g%{Ս��� �����N>6B�3��Hk� g:G���TN1�I!���u�[.�f����<5]����cO�𲏵n~"U������˭A[]���"��/ϳ..{7�k��%@�����O��J�۴c��$PD0�*e��7��<�Q������ŷ �����
�D�������6���wz���i��A����V�hZ�$�mb'h��N���Z7�N�������$�����m��2���p���='����{����6���l5犱���H��R���3��ō�܊I�g��S"���=+ ��RqaD����dѦ�dU��(x�����
b�a]���/00��y�{:iKZ��/�Q⁭>��#�I���gx�sy���p!�K�u����S�TuU:9{��\?�VQ�7P�`��f��?S�$b����-�HdHz�-���nxx�`��ׅ�/��G�Q����ӛ;Q-��s4�M���s�/�q��޹�\4!�@�6�	kv���5DT��hY�KM�֘l���բcs��V��V�I���8Dn�{�ϠN��ә.&S1���2�L�1ݵ�K�yn�`�Sm��s-��I��ȸ�i�3�Z!�@��!��@�3�� ��*��ȞJ�z��Z4�ɹ%z"���xٕ�4Zl�g5BfHo�o�~����"�������4
����|N��� )�o-��t�"���R �I���
�"q|���!���{���B������79[IyL莥8��s��|�[#K��$�����c'��>� CZ�w0@���(��#\�٨��u��D4�%Z�
u>M0��U�>�@{!<Y��ERkOb��U#;��όt[Ό�?�aRX�C�������ÜQ��;�3����-&h��b����)��h�'X��B3r����ϥN�ϼv}YU��>w���A�3��h��g�݃��^y���,ˌH$9>s$�#��P�1.o.Fj�72�9ַ����E��g��t�e�*����R��۽��6*w.ω��*�N0[���e#�'*�Q7T��6A��?�	��h4���W����ML=r�m�?gpD�u�ߏ��7`xm�Z��Lgs�S��-(6�Oq��rg�^�M^����A��j�C�����nަfB͋>�m�k���H�� �kȡa<��?�x���E�
��>��E>��c� =W�%����@>��ڡZX�;@�&�`)�}?D��U��e�R�Tn�(̕ZjƘ���l,.� ��\���՚��l>��^�raV88d��z{B���n��YHuVF�D�%������o����	]V�<[S1�+���[7��\&
�]z�t� IS?�y,hvڑ	&��[ ±�_�Fg�l�$�5۱vT��h�:ԍ��S�y�Y�0�E]!��bU56-��T�3��5v���"	�X'A�l��8�sb%����=RRK����av�>��Ӓ��nêת9�|���v⮠r���[v�$���R�nu�.O�軐��:�
��3�ޯv��[OG���W���bн|qZS��5>H�J��lԪ�|�@���6&h�+d���F�b#B��Z
*��+�9��+��b�19oJ�%n��LwP��ح�*�S�9?�<�L���Մ�"c�>��w,��|������p�NQ�E"r_s���
)��[R���f9�Db<?��QDw�Ѽ�#`}"����+Zݽ,�������$�S�j8K>8u����C�+�:��[��}-��<C¬�0F���8�r�Y<+>A��b�<���Vp���پk!�@G��z�*����E����f!�:KQ�x��R��#��mjaԁ��y3�8��zv�Ĝ:�p�`�d$|�(,���R˰����,M�����q�KP�R��_&�<^X.Ig�E�np�e�J��,���"�t��˕�Hg�vlD2�-?:�J��A�H�p�~t������z�� ��x/u��A4�ӆ�vBuW����o����鳡V�3Q��L�(�m��4K�����mA�=,��m����6W�(W�cM?�к�:��_%� v�c��xh����!�M�"�l,��@�P=Eʂ d>�A��13����>���t�=|���`!��f`;Q��➱j��܀Rԁ��Vn��M�+6�ɱ�Mc�D��Q$�{��6��F��EF�nE6Xj+b�H�yg����Q�1�駃��� I��|�+�}�]k�d���
�f��ۃ:"�%Q�د��#�7˃R:]�"幫/��.�7Rr��{��OO�@�q
���DF�e��779<!!U��k�ț�"PnO�4�ED�#��l���1���?➿_ ���o��VT��::Jb�U��;��d؞9���Ű>C�z.�$W��D�=��p�<�=(��<�Ő�d��%����G��/rR�I�3��_�#���`�� '���|��u� *�(R��e�t7dgL@����5����N���ڤ��&�.�0læy-WU:����HGQ��(>�L�Oc gN!5y4���e�K�Dʩ��S�3T�ԺO�@�2�U��7Պ�`�����S_G��L���C�Td�b-&g�nΨ!`�9��d���P��Q�~k�������-��O��ZA�c�2�I�ŊY�H@��r�&�+���ˢk�r�y�5	z���o|YۍИ�X�z�1���y�չ쑄���܅:��n�s��vI�i�#&�9��)��2���輡#�n�bSCJ��	�럟���Ψ�i�b����@���j��@�+�)ր�nȴ�j�P_�Z�o�{=J".h��r���ZdVgKI#fGo&Q!���S"Τ�"��f`��j��P�?@����""��z��:0Yu��S���6���u���:vj�G��qF(�#Ol�n��\Mo$g���؅Ƴ@\��}��JO��TU�<ž�6A)N�����\���[������Z
@��{�V)�%n�������z���1���ն�/��]���l���kA$�:��r��:����ZU��~�Q��V���Q�X�5�`�Y�@���j�=kKP�݁�p��$��0�ή�!�}�8��j��� �|]Gys���,�ڷ��e�<1	0H�9+���hRG��3�i�V��J5is�y=��ZV֯~�c{��8��k��l��#�����c0���OV'lx[8����ki-��7t�3Q�|LaE|�`����x�t��#p�
�*i����B�C�p�E��
{Fr8<�����Ǡ�N�Ғ��7��'�R���S,�M	�/LR$�U�q�6ݰg������� �,���si'�I�ڝ�[������>���E>"������J�'%��J��� ��ڔk.�ȘWY���X!��"�A�}ӊQ[X�߽%O@�A���T�)Z���'�Cr����q�:F�������r�o����~�F��{��Vk:~��HW/L�f��'c�`}��U��%ȯ��)��f���̓a��"��\�R�$9�R�&�>�c���1O��YaU�Ħy[3�����;s�<����}�2�>�� u�w{Q�H�#�E�;G����
�ڢ!L���KV�
�H�ݚm����ub�9��T��^��В/�cM�?@��n ����Q��pr>��ك7\ ���S�j��/�	�n�]�OM
A��X��ɣ���)��	��L_Î<o�m4+V�������bW���j'�����鲤xV��R;�>�h=�������aQ�?���(������L���\}��ƾ�����iA��gB_����<
��� լ}W�rBJX�ONZ�W#Ă�p��
�ʃoI|��+k��zFdo��>�rW(>�\6`:�]�L�xT1���ٙ0d1Lo	a/Q��A=�R[�����(1��vQ��*����[B���鄣�h���-�_X�k1��;g�&z�sU�]A*h�F��qG"&��s�[=�25����	4{Mr��S�b<�$6���Ws��v���!��d��@�+r����Wi��|Z#���H��ڨC�Q;�Čd�z�P	�o�n�9Z$�v��l|q�b^��=Ax'&���؉��P��K��k#���Ȥst�,�&@��o8m�)Wz(Ѐ ^�!�zspP:���|�Rڄj�M�ӽ�����S������,q*�9ڳhC�ܸMb��������&'ҽ��q�ڋ �?
��쭖���@�4>��U�N'�9:,S�yy�z�	�@|�6��o4���ٙA�p�:��=�"���º��>F�
�R�A��x���vNc�k��s�~�J�9���ׅ����^���]` �-h���Ө|�����x������H�z��Mِ�sB禿#�༵n�z	�
��T"����7S#B�o�����TC��7Ϝ�?��c����ڔ�u.�M� zĢi�y�*		�GNWA>t9.b".Ch�
�FWL�(i�)e� �;r�!���CR��D}��>�� ���5�'���P����C�C�8����#�T��D�(�^蝜P�[u�p��d�bAgO.��b΋��-�0��=遲��͉�ȥ�xʻ֪2�����H��[�d*�#M%P���m�d�/��I�rK�Z�/������c/O���Ԗ��,u�'B^fA]���Ť���?�A�"�����?�^���C��pUC�i�����4Y�ܫ�6�0Mj��N�{���l�g1��:�0���s�F,�J~ۊ��\�;��B���sJ��W3/V�_�i���-.vw�@$����i�l<�����_W~6dF���n���B9D3[����l��4W����$6ݚ�p�1%X'M(e9�5~u'��<��KU��O[�5���e؂J��Co� �}7���/VfN��e�wK$�I0�|�.�o ���EC{���d��z!�}[3s@�Pz��ļ�*����;?H��{z�m��}���]s+{�T����x��ǰ�n��u?�U�Xk���Vgb(uZ�M��y_f�?E	�.m��@���<���s0���'{~B>|0�.YL�4@ �&_�#z����))�4{gg� Z�����6�U��/\R�;Yɭ����Ny�Λ���Ó�lU%5�P�'��&=��/ư�����t2:G�x���Z�}z)<k�.]�Z/z(�4Ôi��Sb���"	O�K�y�<���/��·�!��QՖ�U��	���N���O�Z�A�����������{��v�-��H?e�N�U���0htD5q���]2��CT����*���?�j��� �RJx��+df��Q�]$��i�1�x�n�$�J�d���Y�\�����k�*���aL��OM�)���.�(<�eq�G�2m��,�(I�+66���6�p�3�e_�$"q{.���Z�C�ޡ�-�SK!��L-\��X.�����x�/sb�X�y���K�]��&v�\a�\Va�%]�Hf�ZgX�.~}�\<�C�I'�ǲKF���lF%Px?�W�&�����5�\�/h΀ˣ�{�H��U����c�h�Z��-~1��\�� AQ\�R�LG�W�7�+D�ɱ�� �:z�}��+f�ztǎ/ـ���i���O*�����ʹ�i�fc�K��%x����-3���naV�U�;�?8�W*�t;���2
��f�;�Y���YoR�� ��ج��T��c,R�!�_h��^�a�gaÃ�p�����#�,��6�$�t��ڕ
�4gvb�lF��o����WA��r��t˖C=ͮ<�N�"חκ�h/�u�A��g���UN�̒vD�����]�F�9�#�m�����?[(SH�ɚ��L����m���,Wz��w�6Y��(�GM��"�F>��t�B��cu���:G����Ǐ%���:�PfP?�8�B�y畱���
�3�4_���V����9���c!�0�`�#����5jS���-�!Cjn��xM�W6&v�ϗ ��_�S�8{-��B�^�ݚ�pSn6�8d��H��g�8r�q�1O�N�o"9Zվ�g����]-�]��%�H��]�`"p�D�ځR�e�x���]��~gf�\�B�Ļ�4���ѷ�����	),H�u%��Q�Ri��Ĭ�iH��V�S[5B�;Č�*�?��>[�n�cU����OkI:!lY�P�b���0�O�_1x�{3FS�k"3A�r�_�,�$|*�/E�.��@bHxj!����|
�I�i�SW�;����E�Z
�g�Q:\o�	1���Zҋ��7	7�>8�n�,z�HM�d$�m
q�I��O]��eݺ�|�,���@��h���<Ɇ���⹮�Xm�>{u��>K�J~��ӂ��Կ�.��y/kG��`��	G!�{N ��z2�CM�X�RO%H����o�J�?A��8�9�~r���ɭ:?�	�ǭEJ�r��(+~�����O�[Q:wJ��a��L������q��	��޾������_l�tda3�"������!9A_W&�m	�����v"O�ya��ڦ]�+3n�l��(s;,b�<���v�W:� �����!H��6��;�8���E����L��tPq�V5��H�u>m%��.�}9pw�������^3��ژv��p��rF��
;�pK���ҙ�*16��|�S���P[����'���(��A��q���Y��X�/���Y�塈��cmx9V��>����3��*[���']ѣE(Ӥ܍@V��};�..h;0��v��QS�̣֕�(����ΉQ���}���W6"�hx�Ձ�BY^��P�
��_�9�X}�5�B�D~Og�N��"W��P�Iy
�V�ob�������jd�Ԗ���yW� �\���V��!1
zE�2�d���	��6������T�����E�1Ir�vr�M��#�0Ϗ���0��Ȏ��8���) ���7�tH9�L�Q]:ZU�uv�Y&��H��=NF��q6�	ٷr� �S����]q����.d@�k�¿��@�Rr� %�
�����#X̗͌���sΘ�
��e�ze}P"韙�3sZ}��A,Nq~^�gT=1W&�z�$+���ޤ=�k�� �s�82t���&��)�:8�e`W���y�!�;�s)$��Z���3�4�(M ���<��M���]�;5�q��ڬ�{�*JM��7�f>~�߻'����N�ڄ��?#����|�*�4�M�U�a�'��,,zfy���"|��&��7Z!4Ix�r~s�)s��ȬM�l��L�D$FG:�Ӌ�Rl���1�i�O���d�&s����V��]�@�P�6�P��z�N`١-a��C
���(�^=N�V`A7�ezt���ix�B��#˄ܵH��zb���.݆$����n���B�]���n�T|j��l�ٜF���'�����b���$w �z�i2��*b������A׎�.�O�g���zWeH�i)̈�Y��;럶��q C��DV��7/��9s� ''X�|P� ��pC<�r��\ʕ�Tt��Z^A�P���uS&$�oA@�Ǫ�ݗ���f�D�,���$�3�($���{x���+��ra���U[r�F܍%��Q�&v���\I����s���9*���y�pܩ��b�|^�uu�^_w]�-���<��9أ���"u�ΫT������^{�1C��dp�Ï�j��O�Y)pB�m�0&�1�G�2�����{Ɠ��%�����J7:���U�,��[\��JgZgW��V�W�_�q�����'P�w�M$���A-�l����EϦ_/�dn*�gX>��99}�<��l����M~I�s��*Ѩ'fS�9D7a~�|��<V����������.Wƫ
��ػ���Y w�P�=3vh���be��~$����.VWs 5�	E�<9���&=�|z9�[L����Y��]���⾁F���<�Hp8z��������܏�+�_iԔ�k����ii�̥�2��WX�:��J�|b�7�ƞ�y��Yf��ZE�U".f8C�����Z2�0vs�#��=mY{7;]|	�.RW����@Y�_�w>���)�Y_{ 	v 3�/����.�;U;�����m���X�H5e��ycp���lìa	U^a,7{'C�&�x&/ֹ˰~QK�m��G-c��1�ʓ֩�<�
J]Nē/3�74��(�~��&~	�#�k�E<��/�Ȳ�@27��N��M��&LE	HN�[���ZJ���Ќ�σ2��t�{�nu�fh�ǡI���둶�h�q�h�+5j�Q���0��*s��O%�u�#����DcJq
�+}��;܍���A���?�����'�=���J������\��4�H�E��:���� �l�I��~�S(U�Vq5� 2������I]T�6b�T�,��_��q����EғCXA���@�K��L���OO��1�-/�"EX����Q�K��q�����UAe\o@�%�t�f=d�Xc0}q 5��T�I ���Dϓ�T�%�c�1��)�@��'���G����tV��W�,�c+Aӯ7-6�a"��fQU"	�eA��R�ᚐ{�dױaY���}��8f��.ǧ2ٹ�(�2A�W�-*��Z�S�����f\��K��x�4ϗf�+�t6va�aE��8�R��ʈ�7��k��οl���{f�-S.RF߾�v��Q��m�L�FDR*�_� ^s�g�{�I����J�,��$�}T3tr
t����g/��ldԹh'��~A��*ˋ�tD|j�a��������γ�/�A/��kF��ْb�=�0�nR�?�˳<�;�.q~�pk�(����3V�Ɠ���i/m|��,pŰ����6�,�(:,MZ٫��*�]_�;q�c��@�s���I����Ƈd�ϻP�;j��@��
3@<܁�<����ϸa�նy!�v`։é��
ju�p�;�����nf��M�,u6����[�F{�����?8��a�I��6��t� �H�f�g�L����1��a�����շ�Y�Q]f��D��=���R�")؈����^&�7�]�""@1m/��.H7�o>�V��F�O'n��lY�r[GD�eM/7�eD<�xɉ߾��6oK|pҏb�D�+�����G�C��B2���P�0�pj��V����=�b���_�?�~�V���-Jϰ9�~��Q��ʲ�i��pٕ[=cw��08�ŋd��Rk��&`���y37R���3Du�?I��i���_� /ʟN5� <�R�3��	�dbQ.Rn����u��褒J��BÅ0 �y('
:iW�zpQ��h>��H'��FNg��y/]�!`K��1�ĵ�S���T���������F���70�`r�.��S�2��'�u�~v�d��-!�7n)�2`p����h���BQ����@Z����-��-�$�����d��@{�#�亭��hx�ǒNk'��P�D55���ol���Ye�G���u�F�W °V�&%�Z���nV��s��dL<&6���K2�$�Bp��|�"n-��S����ᢟ��tȉ��i����k5�@�?�
c�̱��&����}�o)d�k��ZEh޹VE!"i p@+��žZ�ӏgrPf9��o��;𱅶"	���0q4���өE#|!b��o>W�t�q�YDk ��II3IT
��|y��!������s�,V{7�x�I
�V���m��#\M�$�UX�@���^�W��5cd0���O�#m���4�uݜ4R����N>��.0߂+U�;��.��!m��L��k�oQ��ު����]X��}8)�rn&X�����F��h~��qr;��6�^������L��[�)Wh���` "rYij����<v-��UB��>ȣ���yձ'��h���� j����ˑ�y��>��s#O��P��_o��Ә)9��T��.�g��p�h����e�롦��瘾A
���J*��k��[�Y�Ӏ�7e��`*DEo7%62mV?�9���I��WG��Oӣ��L�m�x?!
�DL���0;\ШuY�P^ڣ�0L8�u�D}-�>L�������ޭ+r�R�^K���	j�
��ދM��d��o�����_���3� p�"�Rd��e~x�zCEL�x;������ �%�$��Q�Z��c-Zc�;�P�����.��\E�Vņ�e�5(���Z�64�)k�l���Ѣ;�-#����R��۬*6�Ò�8��i��wB^�{�?<Y9!ZF�nd%/hO�Ao�~��'���w�S��Ҳ��[H-\63&�� ��*?���hGΊ	��[��?�����l�"5���v��h�o��}Ʈ���MYP"{���QBp5������}���$�K��ұ'����R<s�2��a=C����Ix�aǧ��u��>���lM�t&��h��`�M��v:��k�v��Ev. c7�a��:���!P�<�"v�O�[��&�')§~"}Ў��qK���gH.�dS���
���s���J�����[�b4���&pw*:�;b_�����bSw�o�Tn�_[w���	dV*b\N��E<X!!�� ���_��/��w=�|�5z�:��5�Qv�#�h��B�)r������^ޕ`�?4ГQ�M9��e[#1<�����+k�,�~��1���p����x�8Fؿ��=�+sV��0}~h�<�L,w	�F:�8���]&�b�M/y)m��M��s�G�J��ʍ��ע�#�c��U�`8Uz�]s��<����C�R��+�w��z�&���1�4pJ�;���z-�P��E���a�~��]�o�Fa���lѹ��t�p4^
薚�$�Ô�;?F�%R+�?�XX=w�.^�m-�A8H���z[��S����m�׮�v������"�L2�
��#:�Ф��қ mG�_28�I?� B>H�G�7S�օ��ȷ>_���z��T��uXP�G���L�F�q���
Z�!��f�RGT�]�jS��%���H����� �!Й8f�0D�r�r���M|������!�������8}���,���ꀙ�:M%+[5d6��/�+�-����'��I��b��RC3��մ��RL6��Ŧ�q��l�?0�Ab�ɟ�3[�t�}�U�Z��ݔ[^�IEU��K�5�@;����ʍJ��O��lka�h�Nנ�-'��H�vw-�V��RΩ9�[?�ڐc�i\d����]�!�(��jG�X>p��}��c8=e�GA���sty[=à~р�p�k��:&ta��n�'$/��d&B�_��ͯoL���̗n`B$˖J������\�{���ǯ�*�~�a�d��*�)�d�p�(<\#q�	e2m��,�Iĭ�6��@6���3�_��Aq{��\�C� ��-dK!]�L-^P���Us�:�/sd�X����/K�N�&x
�\�\V�%]t�f�\3X�p�}���C��I'�ĲK�2���%P:5�W����27�5]��/*Հ͂�{�����ec�j�Z�1-~�w�\�� C�Q\�3�L�"�R�7��D7|��|��:<1}���f��wǎ�wـZ�����!$*2������kfc]K�f�x�g&�/i��6eaVs�;U�8�Y�����bO�2��f�S�Y��ۏR�tQ�����T��TCz�%�R�#�_h��^��ga�V�p�/��L���,�}��$`t��6�
,gv$jlF��o?O���A�a#r�t���=O�<]e�"نκ#8/��DA�m����N�l�v���N�.�F+�##����1�A�(S�[ɚ1�ܦ���zm�7�,W��w��6Y��(�[+M�+��F�:��	�B�cu#��:	����.Ǐg���-	�P?���B��3딮�3�6��:D�����Oz����!�r`������jU ��o6�!��n��[M�YC6&����$�����S�${-{�BnS��\��pU�6�z!�*IHí4g�:@��1Os܃NT�";Yվ�F��Q�]-���ՐH飵]o"p��ڃ3�e%z�/�]؆�"��/'��.s�M7p߸}���M6�O]�3%,��&D���esW�7��h<#�x��V�U���6^�D*���u~�֎sR�Ϲ����O1rVV���|Eb�#�s�fqߞ]��� ^�|���QQ�s�T��]p {=j5�K�R���s��g\UjF��	:��OeR�i�3���='��W�.r��g�<��?� ,�4R�����'d)'��� �w�OJ�b�����I��0��y�ӂ:�����Q:�>�HN��M�g�o�y��;��\�K<��+x;SࣀT�|���x봜��Y�7�c�`� )S!�t�N ����d��p-��\n�c�`�T���P����Q��Q��ke�vH-cί������������ ҈J����O�̎rkΘ��5�PE<���nY��.V��<B7���'I5P�n;O�����<�n�u���6�+�>&�|�k8(2H�������n4�&S�F��E������nMi�����@��+̘� ���ւ����r���.�Z�/�}�k"p��W��P�`Zf?tg�R�f�x�o貧��l�"����4d�E�Php|��S�X
�o���t6�M�`'� ��I�	9
&�b| ��!7Ӈ��V�3Pu7��'IќI���u:��O+#�pk$����G�I�E�t�Xk�ܪ�0�,!рO#�#^�;�u@4{��b\>���0fV�U/���u�!��S(~k��K�����p� �������n׹�#X�ʞ�ۜ��O���e�;C�J���~�g�>u��)n�h���'�vr �X�'���'�BvtqYUit�>�'���~ϱ�����B<���ѸX�,�E��{>�f�#6��PVjgo��ʘ���9eO6�%�+�t��w6����eH;]�7�E�ؽ���*ϪG�ٲ�"��g�pe{ض*�D�7��6��/?�k�EH���W�'�_M���͊L���m!?h�FDs]�72ЏM��%��J;�L�?��ޅ,?���������(l�p^�(��mtj=�w�%�L�Ƅ��ɋ������Kנ> �)֡�ţ��Gx��>ES5�"�;͝^�:�� ��Y%8�����U��ZjZ�;�-͸���B���A�����($��Z ��tl���x�Ҵ�8��-����m�9&��F8�a~�ҹ BQ@���uY�^+FY]%VN~V?o���a��Ɣ�>S������[�n�\]��"�s�f!� �t.?+�rhΨ�	~B[X���f�ڭ���lک@5c,v�ԵhTᛍ�h�ѫ�Yw��o��8�5f>��/h^���R���j��r!����t'����s��DN�=�s�`�p��aβk� �W�O'*�/nw>���p����2�tJ�vA�:�R���'.� ���:fhv�h��ceUv��-[�׈�}�%�����q��{�
'HU� Z��[՝��Vގq;Ѓ�� �pb{�O�M��*AI����Ub�T�o�nVC�w_Զ�0��*i������<=g�l�ĄC�1��kw�X�|���A�:�kQ=��2�%�)��^Z���&$ޜ?�hQ���)h/#���"ߪ+���,�|��8���Wӧ�dh���8���V�{+K'��e}�B6<�gt>��F��8#9�]��{ʔ2�)�YU�T��s�Y�
��4��)���ʏ�`��`_�[�d{��DΤ�
]C�1t첉����m2Y�,�w1%�9p1�乚Oz�>9�|����~+Ǽ]��Fh��SS����l���
O�{�k�Ɣ���F�r�+x-�X��wj2���/Ak�,��e����� �k��oXmS�<��1֠2��ŉ�2��J�6��력asvn\W/b�����oV����W�YTi/�)d;qs����C�`D{|��U7�j��-'�_P�/�ʚ7CBkVȍ0��hhT[Q��+^`�P��u�6��#0 A	|�	PӋ!�El�&��s��Q�n���v xi����7�%����[���GC%/���,�s�Ν�I
~���G�%����2�.��薂i�u;n�^�[J�s5��[����@S�"����Z�����C^��C0�p�ȣ��~1.�b��||>�f�#f�P�*�o�O}��l�9�a��UK
ӤݧZ�	�&ex+ͦg�z�u[�+'�*�2��Jg���vsӗ��e��k*k�7��6�dk?+$��u{�FLW(2���գ�#�L�ĹmQ��?�{}D�K%�g�п����n�z�KL�g�����޵D3�ׯ�
�BO���^"�����jm�8�U.��������#˸������# '�x�����6lFxPE�y\R~a��ngj�] ��=%h_��r��@�EZ���;�����N=��ߟЖ���ܪ�(Tc�Z�D�@@�l�n��ڴ�t��]nj�1��i4R���^8����Z�B5����T=Y�P�F7��%��8�C o*1���~�ļLS�{��I�o[��>\�"R���e �t�?[�Kh�t�	�qu[�O��L+��[l
�15�;:v�
�h�������t�Y��2��b�hڪ5��1�_�]������bW��L���'�Ie�I��s��t��=�U;�>��a��ˠ0[���W�_4]n7/�4��(懶���vq�ׂ�(���i.���s�:��-Ø#�ē��v%��[��È��U�7�E�q�n��I�#H�h�����2eQ��1T޾��г6g�0jFb����}��*q��y�ϝ���b*��o�f�n��w����`��*��j���<O��ۜk2�sV��w��,|F��qáPQm�&��U��)	�I��N�2����P?K�Q�'f�Y~##�oY�RA�+�{,
+��h�ÇͿ�ۤ��8��ن�e+{�B��C�}��<ˑ;n�F|
8Su�]�|,��:�)�g?���s��[A���dO��Yb�����ߐ�C`�6ɒ��)σ����C����%,#?�ߝ��\K�1U�gpa\ٹ��zEE�\�MO=~[_�]1�F�+���������K���'�
+)���$��Q�F�+�G�X	cCw��%�$ҮA�s��^��~O�P{�ӹ*m�X���c�b9Ź�2N@Ƒz�^���(m>�r2˿?QS>ߑ�G���-Ѯ��m�_�:�R�Q
T«#uG��L�1����d�!�l!����~XHTt�~�+S朱~ş�ʮ��,�!�ǋf�����fr	���R�F��?�r�8��������l��ߩ���-���M\�#L}�MK�"f-&�"�G�D��DKb���CJ;�իE�)�৸�Ħ3�կ�h0<K�b�)��J�t�1TF��7��+vb���ܴ�gkl��@R���mJi����ba&*�NN�A-~��wD6`��u�΀��[����'z�c^�ed�*�&��8^1(�K#G��pÐ+�c�?�螒ҵ��t4|�=�(�~���p��Օi���[a7zG�^��0�=��#�X�����K5����D%�&S�/���d{�(v$�gEؾF�J@��i�[ܨ���Hh�õy$S��ɺ�P�o�4���?~����|	�d6Ú�Å�B��g��C�f~ւfc�:/�1�ܯ�P��:��yx�#ˠ��P����I܌V��cN��w��0�M�N	j�Y*�=_�22m-[p���|j��w�&Ov,֩��� �]2≲�+#�D��F�b�� ޴���X�У�B�B���Y���?�j��1���V�����%]EG�^�Y��P�u�^+�� ����3�q4�ǫ�I<Pˉ"P��d��@"%0�L&=3g�K���T�DU��9]yN=a�@  �e]��$�1���u0�{�@����jߎ-��г�'T�h6��nn�Ì4��K�K�����9���c缑�\&9V>x��v�-,��0������3<���ee�ݘN!���-|���xe�����q�!���'� �,N-��3ڵ�`|��n[t�y��I�;���$O J,���u���u~��/�?���7":��(����)�!�+Sdu�/:�XG�I/F�T�O�/��m���g����Qĳ�\�\�&}}��OF�VT�-��B��sr)+��r)�\���	��sR��Wu���F�uW)�qn*����q�z���$�<��ܶ�G����%�IN�����A�q�Eԫ�Q����U%Q�6J��3��������5Ԟ���U�jjL�BK�5��^d��=M`�M0�iY��ڬ�8�j��H�D�X|:a=�\_�.!!��M�?�-�9��	�ʾH����9�R���Pr�il~VUm5f�jh��N�z�7��,.mc#���2rk�l}nD�[�^�0�^�O�#xx�Yj��k���
�Ѓ�|N��EYBm�d�x�����
P�4i�M<��*����)Elґ
�|�UB^a�\����{�/kt7-.��/��4?,��M����$�/Gq0P�*��u����,(K��0/���֝��'��e��yO��j>�����g�J�8��&s���4S�wH�kk���4h#�-C�Ϥ��G��TX���%�\��UR��6s�q���\].�rY �����:�#4-����r"���^D~�F�M��ᑟ:E���E^L��뤃�}��KY��$���k�s��wa��B"���o�_9e�W&h7��J�n9�O/ďa2����D$3�r��1H;Џ$<���5��{5� R3�I
H7�)��g;yʑ��vÍwq�L�t|�4�VY0H��AmIcp���B9�!�Vzу"	��Xڼ�l�����ﮔRpo���v�Nؿ�j�S'��LU��[^��LU�LC�AGӥ���ɀIn�|�?�&f�	"��&,m1�&V��ַ�j���:��򎛱s3K���� ȣV.?H;��Hh���2�q���~Qw�c�z
(��R�rlr�7�5}i�ž{Ɖ��ե�B��o��R�
:���]�\}4�&BǸ�O�rN��GW���m�
Bo���}��d�1-����W�6\3d^�����1���VT�dNV�	}y�:Go��ξ5�d��1��v�8G�q�G~�sm��x���o��9H�ܝ��-?���[ce�E=�p`�]ޔp��N��&����W=r�I��H	13�r���S��I�A�e�Ҵ䶏#����@ܐkr}#	�.�%�e�#|}c�;S��ܿ���ĉ���PF$�K�%Z�����D'q�>^L9�=>7&AEP�HJa�r
��ȵok@�,�5sln�tݘc&�+M�?8J�W�J5�д!�0Wsͽh�~�xŹ�Y�X� M������;�5��6��2�q'c��P�˻NRM?6�,[�
�p��'sYM��� �(�H?G�_슄�N�"4[ZVU�*'HΕ,P�Gy���FY��[F�4�Oٖ9�͜��
������0Úh�Fk
��/~R����P��s��N�sl��'�������ł�t�����`���-�S��G�i��������[��zK;ٍ�B��@#�h���z�Ň�..�H�i��({	��BD'��uT V���6���� !P�Q����o�:* �e�i�B�*����dA�k6.������W�%i��}�[;�̜��2�C��Dz�'��H�]&BuM'|�eP<���vC�Ad�����^FT9���_^e	[P*��uw�����QAd1 �'�܋�eu
�M�P����+��Ly��%�sx�J�������%1�[C*���%������,¼I(.������॒ VjL���� 8u�^J	�Q�:ѢH� �$�^ �"� <��9�����^HC�Ap2tA������uYMm8��q0J����|׼��<�D�Ʒ4׸�B���	J�?��m;+���VJ���WP~VV��_'������˲w0i'$����e=�lYe�ix_��)dC�a�f�H���f�3���������L��V��TY� �"tЌ~o
1S�Pm.��q�9��GY�Y�t �	e'+�,ڪ$��3�>4~z��]A���	�24	���@6�-��w�3�"�ߪx�2-TD�OM�Nё|@C:e�{��|�1H�F����{��^��gҬ[ߢD��d�@�;�,h��Ě!��W0#��aOK�l���$�b�Б���(�9jmx�I�A�]�\]%�����݄���eM44N5䐯�ǵ�7�,vٓb��w�ލ�����NA��3nU�`�)W0���V�I%����� �������!�u�[��*ɨS��ˡQ:�L�.
B=vY㿚�u�i�:��G�XFyF�O�;[�i��Yg`�t�_̳Q-�\��i}�OZ�T���폖�b�)?ɀ�N�\���� ����ô��g#���)�B�n��;����zMn78^��o��<��.,��]��|�gU�4���)Hi�L��U9��5��G�&'�55h4���Y��j`�yKPu��r�M�����a"׮�B1���/8�C1j�/��؅#|NgZ�%�B���}៷S�Ǽ��	��Hh଑�R!�	�d!ri ��Vi1J5�2|���$�K8r����c7����kPl��X�!_�R0��vOg��x����ɿkڀ��*�l��D�|ⵐEm�}��9x"ل�tZ
d��iK���󿡳P�E��P
��hiAL�BJp�h�V��C��7����C�&��,2�uMZ#6�&$d�qD���8
��w纫��,<���Ė9���2�x!���v5皬����>3�\����J6t�:��w�u��-Zk�;��H�e�����3n��A:���Xy�c% ���j1��H�:�a�@��]rmX�с:�:����,���;r��U�~V�q�aׄu (:/�W��DL���8<�������x?��Z�j�����y"aהH"��c��� 9�&|�Rg/&�B�O��aF_��� 3&n��R�;��<Nqa�.��� f}���WHK�-��;�&��7UA��"2LcH�{KV�8�H��Um����"�9(T��j�䃡I���a�P����|�*͒��p��E�Sl�~��S����`�c�F��$B��A[ )�)�ɔq�ۚ�:�!���P���)m���V���[�����hK����Nߋ���-���J�VB�;���h�Qk��dK��#�Q�Z����(f����s�˚K}}���@�  ��9�!B���>}�
NKM���}H�B[�O�%No�WW�� �{>
VR9o�[�c����Cd�쏅�ݕW�}\�6�6��I�1�{O��PGdb�\	����N��Փ))�I�$d(�1��v*�;��r��CC��K�ƾ��У�������p�t�F��|� ���/�]�5�Ȅ�b�&��| �A=5u�)��	�U�r�4XS�%g�Sw��Z��b�#�*�կ]   "   Ĵ���	��Z�Zvi�
X���SeB}"�'*<ac�ʄ��i�*b�P��?Y##��V�x�ƀ,F�q���9�VD}�ulڢ��<�2�Rl��#��)w�,���-3ϲ��pӌ��=	��/�!6�_��򵮙Q�-�f���U�	�l�4���i�j˓r��k��k�,ʓY�8%�5{�l9��#ДT��hJ�GVj7��ǟL̓~��y�hl݉뵐�T�EM*;�h�����c���H�W�ʥ+��O�I��E�y2� it��TF�聓`	.��k"<	v�?�d��6��1��C=gv���a�]t��O�4���D��EPF�1b��,5씑�#J"�jFx���r�'�v��'�j�8�+Q������AO��A��+;WqO�<f冿k��抗9��(�i<� Gx�Gj�'�`K5�U��U�B��!Nȸ�Y��'�n�Gx��r~R�\�1�~�BV��]��1���F��O��P�r��#`�������)	^��"����:�ExB�X�'��]��6u���ħ� 0�&k�=DzNb����ች9!�'�hY�dL�U���Iǅ�O�D��'��PEx��e�'���ɖ�:�V��C���r�Q����	%��o�F�'��u�;�yG�(-Ю���@@>����Z��'�Gx�~�dו��$��i$(�)��U�J<Z��'C��Dx�`�@�'�l�9U(��j���HB��:v��
�'8�W   ��$0�A���y�s@���W�����`&=�T���P\'X�Z(^��z�Oy%�#P ��k��b�s�����t�Ι�L�j�ޝ�Fg��m��n[Y�� }��#}�h�p�9ͼ����F��{�)�7�t���X�.ś����ߴ��(ҲJi��Pb25\%P��\���B��������:1�؞�Nף.�Έ�wlN /.�j���
�:[�H�Pz��k�a��ħzH��P�>N0\�ߎ�W����[E�"��8ZL��?<S ��Ce-������W���O�Q��N^�ښ������{�����`<R���@d-Ű��Р��p����[��.#x����^���GR��5YY��!^�B;�Z�#T�og�������TO	*�GuI�6�1�镗{[�3�`��&S>��r���EoD���B��upݷ=�U��CK�R!z ]6e����O��ϵ@R��z�C~�!�鎑Px]@E�T�0�MN   >    :IZ@-�nkZ��&C�'ll\�0�Oz+��AI��e���X�'M�X   ��Jn���������-�q��   9   Ĵ���	��Z[V	�&��SeB}"�ײK*<ac�ʄ��i�*b�\x��d���R�`���1)B�[c����#���oZ��M�q�i.L��$�>v�f�*B�A-D��0S��ھO�HL�'�֗�M3��D��Oz(ݴk�@���M#_ޥ��:~��E�'�ha�$C�Ʀ�/Of�ZR�[&]ȝs/O$m����۠�AR�Z=*��)��$C'k"DP�MJ�?��']BWA��+r)?a"��>��Ac���0e���WUN����&���"<ɡcm�`��j! ����:N�d N*�䄺�O,��H>1I�ZdA����,�
��D`�<)��)�f�J#<��l� Q8 ��@K�^B��� `]' q�P����?
b�I�S]�0�g�G���ۅ@еg7��'�z�Dxb)�P�_M���ع"�����&#�pmZ�������IY�Z�ePU��P��'�Hu��%�IRb������8�%��	^���eh�5K����2�<��G(�z������(dH�,@2o�1?��(�욱}���0F�I9����N
=Jш٠@�|(o���1O(���������$L�3�K�� �ED�N�P��_�#<9� 4�@u?�`�H�g�V9�2��x�Y#����
xt���O�ãH��Mk�4��	��Z���?��u�?zn>�����&��4�_~ҡ�j=��Dy"�	w���(%p\�(Pb_Y`=���K�N����<ӧ�I? ���R�	�X5��!�X�vB�ɾ���  ���[�JL���T�}�L)A�K�Tx� I�O֭$��:P��	eR"0g {=����O���O^ʓ�?y�}R앳����b�,>n\�$`U��=��|2��\K|Dх�X�zYh�A��ޠ��'�a�ܸ'\P!���^��� ��`@v���Y 
v���>�Յa�rAэy"����
�t�2�  t���B�����ȓ/�F �����?���,=�8��G2LO���P-��W_01�ᧅV��7,+D���W�b�4���a�%y侅b�f%�I!�HO�ӡ���u�ofi���<@�<�E{����b����?��@�h�L�����%ҷ�(�I6t�%ڗ��|�-]*z�����Aɓ�r�͹�y2B[IVB��쑤C5����MH���'4ўb>ɘ�`��
�����O�!ז��#D�������.�L�y�ϴ("��qQH?D�<H�   >    :IZ@-�nkZ��&C�'ll\�0�Oz+��AI��e���X�'M�X   ��
�*=��'�8�Xi�#o�   		  �  �  f   �(   �pA�����Zv)C�'ll\�0BLz+���4��'(yc�F'���) i8�����j �3D	�@��p�^ *C �����&A�iέ;#�<1æ4Pv����$��	�h]��͐�*�{�/R�3��:w��O>�9�d�O��;�Ɍv� �B?{�x򗭀N����dRT�Ɂ!���S�O�l���h㞐z��E����=!�c��%��dD�.j"bT�1cD�J �V���	��@�*�I�}Ϩ���(jp팁.�t�ES�@J1q�!�$S�e��Y�CKQ:{�>B�./owazr����7D���P�~ȴP�d-�Z}!�DƉ�j���˪YĚ|B�,�/OH�O�Ezʟ,���'�\�bi�R��#��x �g	j�'�pd�9�ɇv���
t|܈3�݃�J��)]M�bc��@�FD�);q��'�"@3�ӢXQZm[g��?�,T�	�'�J�Ȱ
��
f!`�H�:@��{�y��)��
2J�%�-�s����/�B�VB� b�\�S��
l�<���R�+�p0GzR_>�؍���:xƐ|BF	�- b��a�R5�?����k1OT�h��S�?���3a�'�����_|0��H�J��)Qk���6�� $4aW��*r!��V�|5b�I�(X&ܢ��4��H��I P=�Ȓ���=mL�ԡ#"�C�I>#R�	�M q��	P��ɛY�����f}�3�|��'ˌ}3t�Ζ n~dPVD0x�Ԙ���XC\
�'�C#�@!3}r&�*VȄ�ur�j3��ÔGn���KL�g�}�N�;q3^	A�K-y�d�oM�6%��t��#&�}R�_�!"C�oYfd�� M�bT���?����?�,O6��4�	_|���5�ܼ-��[��]�"@<���D�JF�!���ޮچXS��VX��	q��D�=�O�){a�Ă�'��a��L���ţC?��	�����$<��!xW���Q )޴OF�9�$�W$b�d�Җ"Or�f�!v[�� A�5��T�'��O.�6"W7%��<�V�܍?�"h"O,� 1%���y �(�9�y�P�$ZW����Q'#g.��2.٣���Q�	��I֔�<�`KڜJ����J��n��TA@��s�A7H�z���q��%NL��N�zMq��٥O��B��L9��X�&�fI���xr���6O�O��>�Q��%3�#��E^��qa�xr��?����䧲ħ)���iWlV�v�����CG����=��Ұ<)qhUq<����5u�P� �(dFz�՟�}���	�fHA��S����`A G�L6͇��?q*O.���@ӽ����%œ cf��m� �^-�GI�:Qq���=}�k�ǰ<�F��#nI4����_ɢ��d�^��쉄�3"sҥ���U�p���`�$Sk�83�y����?�}&�� kכEu��"*Q�>�z��(D�井aɖ9���W���O�lXS��O:�����Gx�'T��'�0�6���&q¡��t �����4����i�O����O.�d)�.�L�O��ĐO�4{�+��DL pp�ͦr���P�A(%��~"O�
.�!s����o��	e�)�D�$d�}�S�`���0=�Q$>G�]��&��fE��ғn� �I⟀CH<���?��}����8G^�B��Â^�|=ȷ�ݭ��O�q�[��qJ~r�@�:���K��;�Q�E�&w��'�����'��	�]z�' ��n���"=!
(��ej�
�.Q	���?A`@Z9z�������&Q��:f(��D/h��x0�΍@G@%�"
�~~ay�� �j�U܅���$T��X1e�T+E,��Ȇ	RoayB�R��?!7�ixJ7Mr��Qɐɂ%`�"��Mu~��cp]Ty��'U�O�DQ��߸! �#�I�S��e����LM���i��z���a@�`���MʏJ���`%8O�O��rj��i/1�J��O3ڑ��C� ^��+�;?����D��@�ep��L>)�̞-.��m��&N5B�b�<�`֨S����b�:5M��Y6AG^̓�hO1�LQ�'�tl�0.�:�;q"O���(N(x��QL�7-�tm�w/$���L��Ьy2̊�zM#�bI*]�d���-%<Re��y�������Ђ� @�#��C͘�:��T�Z����k�>c����0h=�� �D�,���%c*t|!��.d��X��)�� ��������ID"�Z��]�0!Z}�dĶ+��B�ɴ/���P�W�Xu*�灺B1��D�T}��(�V`�'����-�q�~���D�k^u��'	�lذؘ'�P9�/��`�H��4 �?��� ��H#6y��Hf2 
�.����b�fYJ��ȓZz��@���mcV�S�
�9D$��
�'���!�&���*����8�~�c�<��'�rP��'��h*r��Jw�����'ғXvm��'dvdR��č���2�.սw�e�J�P�$�X* �Rc�<C��/�I�������J]�@�a�5 !�D�WZiyE��Hl��9a��2azB��ذ+\� �,^�V����q�Zj�!�d�6]�ry�1�S3_��T�em��&��O�Gzʟd,����0���Ɇ%U5Xnq���K�'U|�+��2�	�-R���_�g����S �Q�DK�$
�@/�b�t��i!	�q��'o2����s9,r�����9�'*+��A�%�L��ۊ�~��y2�)��l�$��ƃ@�& �1�g�{>�B�IH��x�J�O�b=!�]l��Fz�]>�j�r,�E|�@���6z�B�8`�-�?�P�;v�1OZ$�r�Sv���m�x���n	��P�꓍(<���ƝT�y���b���`\�
�!�$�+M4up�|��93#�S�����I &�D�{a�U��<a��x�B�I�citH���5U2��`��D�j���@f}��9�8��'aTH������(�iU�]>�Hq��'���&���'��5h�f�/���4}�.XS��xPd�����-��-8�H�5�-r@�1P��{X  �ȓW�pӱ�àH�ܩ��X�6�j���'��bMP9> �(�Bͪ4��Ĩߓx��'l2��l1"Ⱦ0`g	
P���k���2ғn�4�2�'Cܕ
�d��7?L]YaJ��F��T:M����"�Sb��$�/�IX�^�����C��6Lcq�ʈq�!��߄)i�V �N(��c,4������'�Z�ҳ�Zx`���œ9�>�j�'��cM�)w�]��/+'�0)���?�S��.�.I�:���B�n���H�)�9+��"=A�H&�1O~0"A�O-��@L�$IT���^�N\��"��$�������L>��qkH�J��[ Se^�p a�L�<I ���$�`]I�I՛7�`�4FF��hO1��4���CzO�#eD��̰��"O4�i3m��,�b6��&kҠ�h(ғ��)�V�JvHA#�F�Xb�]�u�"����	=Q}��p�y�I��x�*�O�*=���I[�h.P��-ɇQq�+��';����B�q�}��Ą�p��DY�'1��k��O��|a��딦<L�\����&<O*ɛ&�O�p�@�kE�3X��5"OBܟl�sM���zG���D�$�@m}2�9ғA��'V}BC���/��i����#2ƭ��'>��s���ʘ'lE�v��m������*t�jt�n��]� ���N��I��^�Np<�0#�%�f�ȓF�X����� O��&@`�@�'j$��C
'-ft����*�h�:	ߓB��'>X��D�=[�L9ă� O�H�����:�*�li7�'9��#cI��6;�`"c$ԲS�p��O�xR�W(r^b����g-�I�;_X8jG�^iޔ�%��:}�!���pozt%�4�����!ۃ xaz��d�OF��9BE��'j�53��qN!�$]�p�)ԢNg�U�I� Q7�Ol�Fzʟ$�g@E�<�;���w��x؄Dx�'B�;��6��D�.O�y�z�y���Qh��YV��=cHb� 02$��Cq�ɧ� B�  �(��b�J.x%�5"O>(��f�l��P�!$܅X)�:��+�ŞF�����Ȫ�Ȁ�Q։?��Յ��.i@6�)c<U�#]��60J��d�|Ҥ��{�\#� �v����'��L�l���c���!=§:&���@a[� @���5J��	��Q#
�z��	�vօ�ćZ���)#�B۫R7�C�ɿ]��@��A��X'��y���KF�#<�ϓ5e�<(w�&n��j��D�j��܇ȓk�.%� �c D�Bwo|����	����j�'��O�]9���%��-��Cٔ1%r�І�O�M࢈b51O>Y����L��'36!(5J�%�<�[�bW�:��?D���'�ϑi8�xR�Y")��%"E-D�h��?����Q얷.|�E��bh<1 ĺcHf�kŬ��=�l� M����M>�C,��]۵X�-&��aN�R��x�������]-�?�5��-gB��Q�)����y�Ā�Q�dЎ�X}*����Oj��h%F_�bf\]� �=U[4 ��'{�$A�#��k��9e�n��ӓ��'}f�h߇s���	�O	�ag��	�'�ehq#�
=��

)a\�(���$�S��j`	�H�fDǺ:}�84fȃ+&�"=���{�1O1��O�^��E�џ����cˍQ������dƬ2�� k��L>	���;F�X%쎠\�6yѡ�u�<�T�~�Z9+��ޜs|6ܒ5�^n̓�hO1�A�!ŧI���D��&N���g"O��H� ӯAh� n->���bL:ғ��	�_��Pi��Ŏ����LL|t�	\.���y�6��f8a���M8T���*iD^t�F�R�
Mk��'��%B�վ,f&DR�Prw�B�'h>�B"]2���+��L�l�0�q���!<ONȠ�ˀ�FyR�1���--ڜp`"OΈЁ�ݍZb�� u"߅yp,��@�'�:�RN���HI>��f��FJ	P�۹+��6��`?�t+�;=#0��<i�/=s�%�\"G�X�l$�('kL�.�XqKF);D��ZEJ�r��	���&a{89[�"4D��+Q�b�1�m����T^Uh<Y2�.✪���'�|�A�s��cL>	�
�/�h���E�<pâ�س-Cn��6����C�?�F��P�THQF�B+  �E�S���N�<T���d,#��O�U��MŜM����بq4Dt
�'�n��V�Z�r�0���/S�u~��ӓ��'6J���/ʅuq��Ң 's~ �'�i���GD��Ac޶L� �k��o!�S�H�%z����p��8 �7
~�D"=�͂+�1O rG�O��};w�I�RQ~1���Q�.�r���E|%���L>q6�� �p%+5Ř*bꌳ3BP�<y�M�B�l���l�����ȉ�<y����B��+;j�msg���k!�D�p�VA�$β!�T�dյ9�J"=I(�xx�?��L؝$dR���h8!��9� ���T�Ɋ�Ø'F�d���˧���Z�����č�6�Ǣ� 0%�O1.����Y�M(2x4N[�\��
Qd���y�i��y-�xb�P:)*�Q�P�ˮ�O���D	Vo @2(<\/
<Zԅ\� �!���ZjJaa�d��5}ܤ)�$
c��>Q��I���v��[����kTdM:��S�zq<��B7��YՄ~�R��aX�`�\�4_��@��?�L��D�M�
B䉉}��p�)�P���	��+G�C��:&m>�P�3)���wGG-)���*@|(S��YDN���f[4%le���1��$%�� k�%N�~싢H��6��?���	dd���2��uK�(�-~�쥢�䇱'�H�Oθ2Gj	�9~1O�4��Ԍ��(J�,R�I�m� ����y
� �%$�Dy�hz�E�~xd���'��O��R.V -V����C�}���"O4�`BNT�oS���Ќʺp"d�#�d�C������F�Ɖ��)X�#kRM�@
b`��Fzr�,�b�$�r ���s3f9yV���oT8P�xy�L"�ɋvP�y8���|��	�f�5fY o������O3�yRkеC�A�qǇ�]T��0�fߝ�'�ўb>A��i��H��Ք f�*p�9D� �F�[��"�w�Τja��;S�[�'��S��'�F��ׁ��(V~	�#m���H�k.��r���X4>���BM�#�4��%�R���@l�K!�u��l3�O���P���u��� 7m��8�\�0�"O��eA&/�D�QkD�w�ļYP��Tx��ƍϩ8�`���RJ�X����"D�P�ƅU�[䈍Be�N*k>�!�c�O���'ö#=�3�|Z�)N]���UM�Se����':���go��'H��e�܏����5#A/��Y�4%����&y���ȓO�D��Ȫd��U�$E���7���̛��-�hD&�~@{�'�8l�I���e/}J���b��'G&�c�Ȏ0�$H�,Ÿ9���[�R�0ғ
�t���'��iP$)�%LJQy���FEƌN�	�d§4�@b�����%����Z��C�)�?uԝ1�g	
�!�$��~hzQ� �P
� aF�f�az�dUE�J��h�1�:�:ƅ�k�!�^+)����BBν� �2u� �T=�O8HGzʟ*�)H�3i��	1eりO��i9���E�'\J���!&�I�+�n�I�)��ـ��5] &u�0ɗ
Jjb��� ��T�q��'��)PС?&��������%�'�l!C%�	v�q;W	>dк�yR�)�S�g��E�VZ�\�k��(0��B�ɸB�$�釭Y�g�5k@���|��,Fz�S>5��b��?�J���=�� 4FQ��?-QZ����y�#���`��&�LN4:笕���Z0O�1��4� �'���(u�N�M�̩���y��8�'���A.�e=��Ɛ�m�حˌ��#<Or��W�{��X��%�H\ �"O��+�k�D��hS��
!*��'���#�� jH>�f ���Aba�J�{�,����y?�d(К�, �<9F!ԇ�zT%��BWO��"f��*Y?��C�#;D�8�3n@ }�Rm��*A'H|���9D��bv�J���Q �ݬPdF<{�kh<���ݫU<r-AA�ɹ+`n(��QW��(�H>ys(�a�"�`�)J��^��V��i�����)�?Q��	���q���0H�u����P�D�>s����ăh\�O�l�Hw!�E�>�k�B9Z���j	�'��uFS()vLӭ̎{��aӓ��'̪��D�l��$��O����'E���ԡP�|tf�U��Cm�ቊ�K:�S����`2t9R!�80�F��G�s@�#=9W�ۏfE1O1���O
8L;��-մ��cA2��*��d��+�dÉ�L>� � 5�(�s4�N���% v�<	���2�lH㱊�>� ��k}̓�hO1�hu
0�
� ��͸SlY� ��y�"O.)9fbOI(bx0F)�/鸢�3ғ����K��}"�.%.�Ht���y!�DzM�O�}�q�o���D�DV?�(�2J��qQ���B���#����?����s�P��7��"ۘ �!�F�<1�E��l��.,�}s%ې�x�Fx��'9����Y�j���FR�$p�'k$��R�߮_v�5zGFC�ϺM���l�	��HO�e$�L�k�1ed:A�I�4����X�f/�}��c�H9�-6E`��O|���aC��	qƬ�z���ҥ"O��4o+/����kY�(�Z	@�"O� ��93�X/&�ælb�2�Yn.4��#&Ôe��p�8�0Q�D�8|O0�$���F�.�=������$���#��%�HO��3H���<�$MR�)����H��J��CĎ=}҆L� ��`ʋy�O���R_�Ƞnè��P`	Lm�}��q�D��$��d!`	PD�.��h���e�~�0�(�
�&Ї�;��ȓ776 ���3Q�
5*��Eȼ��?Aq�)Z� E ��D��m��4a�2I���`9s�_ ��'��������3�ͅ.g�� s�[�Nn�@��yB��,n�$�}&��
D#�Q
����A�2}� ��;D�(�W��)*�x���&��<�v�+�N���O���h��^l�KS�H��"��'�0Ly���X�����/FCP���	x��7�Ia0z����c�����B�p�=l����'�(,Kb/Z"�Or�87/�*J���B�©=�И�O�kbH������ ���f�*H�%$ye�g�ɐ6��|�2�/Sy� ��!;����%b"UC��'�~����6�3�D�9Gy��PD��/E�2�bq���c��P�	B~����?ͧ�HO� �ud��=!����(�b1J�"OR��T	&v�6�/M>$ r��O����Dx��b�b_��r��+��]��$^����`V`ҭ*n�l�}�'��M�T���I,���bSbs_0d��d�x���Z1��1��0v�>&�d�牥6KZ��*�E�(���h�v���1񃘛~��iY�/N#?�zd��I2�m
2��S3H�S��q�����O:��"���'d�0��5��ɢ��R.] dq#ߓ1&�'b��Y7�I(R]���#:��Y�{rl$x�\�0��`S19�h���{���Zz�g�YQ2���p�\��?��_�0��5�͘�?y�O
�A1�^�nT�� ��p��{��D�$'t�Z�ЙJ�~�$�<,O�Tk&�ݺ#��}j"�E�<�d��PO�%D �_��3`�wX�Spo�O��$�>��E�����2fL;U����e��_�հ=Iê�� i����^ V�1��X�b���)2|�1��E���AW�%��&�H�?!�{��2f��c>a�H����r���ur }Y$I��N�^ �A!�ɴWM� ����|�.V&C�����<�v�1�댉�yb�P(��ۊNA�0�M����y�)����P����= ��`�C�mv�B䉈 ��1���Z�M
�$���/uPuFz�U>)ҍr�~w�P��'��\	��?�Rㅿ�1O0�� �A�m�C��ɦm��/B)=�D9p�Ŧ_�����TWȜ������Ĝ'gh!��.Lu	C"�;>�����K�W_���牀j2�X��6v�Y�1�3^�B�	j8�;ç�-OhΥh7`ך�d�p}BA#ғsp�'���E��LC�QO�(O�	A�'3Je��G�2��'�����҅��pI�p�ǟ	4����]?e����S{�x�Wh[�4��]�,M>��ȓC����'@ta�%#���Y�l��'�J��r��H��ı7Y*�Y
���'�F-Ó̋�|�\�Z��W�4]a��4ғGʠ��'�6\jq�@)%��EȦ�[�r�VD#I�6k�kU~c�X34�,�IQ^>�amǽPU��t��-+D!�D٫o�H�	!�Ѩ=�ұ��@az��Dƭ~� y'�I�s�t��4���H9!�X�]m�0��B�(�����`�O&�Fzʟ �(A��4ؒ�	fNZ/'^a��f�'ڬhۇ�5�I{�@�)Ŕ"�� &�L�;ǂr�c�\�" Ȃ;q��'ڲ��bE�X��MP�+"� k	�'��UP5J��rN���#�te(�y��)�?g��I�"]�/ز��Μ�
�B�	��8�T��N�rh��-�yB:�Fz^>:�Rh ^���`l��?��'�P�y��'S�u� ��   J   Ĵ���	��Z([F)�]��SeB}"�ײK*<ac�ʄ��i�(b�Dx��`�p�m�Z6�$���CA(`��Z:eN���4Eӛ�p����	5H,���J�ȕ���"`A�(�*�:'�f(5�I������iq�Q�g � x�t��6c����OF�Se�Ֆ�M��W�d떯+!�Hqc�]�����E��f�����\�VaS�)���An	��M�O:�p��� �u7�vyu����|���b��i+"�@$)�&(��`�=i��,;m�	�@�LzP�!YL`8S��9OO�a���$^���	$���!Ȟ*�l����L�4�bb~#<aB�3L��* -L�E�B�:e �JE�ɻSV�hz�U����5)�D72��1�"}�Ii�'5|��=a � �kC� ��*Y�`�Q��-\���C���;|���{w���S{^5�'�><��`p���(c��O����$<��䀢]�L�p�j�Rt�}i����<��	�y��ā����Z�6� i�jc����P�zv�X��Ў�O "��q�,�ꊌ �z�k�A	�<���&�,O")!�Dku
d-�/y4�y4�O!����ģ��]r~��ɈR
�)����BnH����B?"�N��BO�=ds�Ą&*�~Ȋ��ݦM�O�P���p�ɂu�6���̑(0U�a���7�˓Q	|�*A��\�GEV�3�I"� �S,�E:%h�f9���_Uf�	A������I�|�����Zxq���O�B��C�I�36�  �����:�0�n_�	� \x!a��&�s���I�C�d�V	D_@��˄��%t8��J#}����{_�y��ӹ���(�@A�p���
CЁ͘'�vl��'��`�0#���s�M�?F>���������=����'���'~�[�lרOt���r��qA"Oh�#�UM'Ĺ�6f�?j��M�C��y��� �O��E�O�f�Tp���J8*9�2D��"�V�j�(ԮR4|����ܷ/���sO�(sv�̝%�R�[����tCLE"AX�C�	����aː�7&f`�BH%8�H��3����N+Z[^<���e���q���rUR��!��Q���
?.�I!�(#U�Y���!\O�$�=2�^��� ��B1�) ��@�I'=p,$�����&?�n4�'Z�����;J�@�c�g����X�/O�Y��Ѻ@�   >    :IZ@-�nkZ��&C�'ll\�0�Oz+��AI��e���X�'M�X   ��i*dJ�M�C|\)2�   /	  �  U  �  �&   �pA���d�Zv)C�'ll\�0BLz+��[�)�o�g)L�RY���B�	+� �4��Dh͙?���ₒ8#k����X�"I���T�#m2p�(�ob��Q"T�Z������&3�bx� $�aJ {Sɖ �$�y#�'Y2�|b�'Kr�$��;x�Ç@��
���!b�{��*�d�}y^�[4G�&k>n����UaqO�=�!��O���𒇊'�bŌ�1�݉ hՍ�Ѹ�lX�G9tb�8:��'�i_�8�t|a%ȚS(ƀt�׸& !�d]�����G	><z��/Y�azr�Dۺ����/��N0� �/M�!��5�t����gA��{��[0-5�O�=Gzʟ�����B+V��,��%ȦZy�i�6ړS0�K'�$^����� ��`W�ǿkA�g�{1O�E�f�����-L�D�۰z!���0N��@�Ň���)�N?$�t��))a��l�<y�����,�̍��B� ,!�nQ�%n!���GC0�a� "B��RA�Ͼ�t�=�O��O�un�?�6�q���}��JP8O��
t�<�	e�V"|��-\�X@&�B7��='�Xj�fV4E���F�d��p�f�i�������#NPY�0D��:/�6uZ�r�D���p@SC.���<Qq��=vH�Q/^�0��ݠ ��}�<������8HD'ڄˮe`�"V�<��O.PGz2�2���m9T���W�]�B ��݊���@p	�?	�g	6�"ܤOĘ9N�u�����P<�N\�e�_54�\�I	 �O�`�E�Ym�L�
�Ƃ�?�\���kT�lVt���+:�Op�)v���j�.D{U<@�s��T1"�2�'��'*�	��,�>�SH�2gB��h�HD
6����U���iO>i#V�_ȝەAT�C{���6��E�BHa���'��q��N���kR�F���ÛA�RLC��>�#�b��C�y�`ڛ��'�L�Q� ]$m�Pl��],a�6��B�BK���\�p�¶�Ӿ?�&��	n�� x��v�X|0:����N�����t5+���u$�ir�ǜ�
S���?G�)*�G��R�LhT�G�L�p鋍{b�אP����C��þ����у*�"��B���l����;I�v���ۙ�q�Ni�O<ys�Q�`��~m���x�E�u�O����P�%G�5�^���J�e<eʧ�x��
�?���䧋�' Т���~����&�� =(�L�=����<1�똼X�Y�������Cl՚�HO���)���|ڤ�΂&�Yju�6@p�؛7�^�[p�'��I9{Y>U��4��'Al�qH�S�hG��zFFI�3@_�S� �K���W�,,O )�"GX�rI�E��#�(F�lH�$�d8-6ayO�2b��=�POO8C?�� ��}�)'�����Oq��'
@�RV˓�u�<Ԃs��f�����'�Ұʴ�2x���r�_�260x������a���)��	�|^pꡃ�*�FU{���7%�^@�GӹA���'�r�'��	(w����?�%㝟b� @�M�1�=jc�P�&tpU��\��X#��ןM�L��'P*���o�zd�M��#D=y�T@C�?LO$���+�@�z�KۖK���
0�G���'��O����OXc�t9W���B���͍�S	r<�AF;��t��'���v�@��N��LIC,�/;�zM��kL�	4Nzi�I]y"UE� k��'v����e,��b���n=V`)2�Q�?�t�$�<9Q([,�?њO��Y�&!�*x�O��*��N�/��1dC��bC��8��'ά�0�H�F���O8��@��
��eѶ!����'(�9��BB�&��\7mC�"\��D$P�p���&Ο1�6Е'����iC�S�`��&j�?S�*i�c����D{�O���j����K�$�'H�-T�X �FI?�)O��x�C�,��d�O~�'2��i�~�	UBq<e���
4�B�YWM�O���2X�`�@��u����|&�l�a�SO��0�θo9�+�N=�$��@�2�(�A�<p�'`���N܂"�͑�� ��=9Dp,�w�x2�I��?�MU�O��O��8k�.�9z3> �6H�4D3 �؍{�'�ay��^�KlU+��Q|����H%V��UFy�=O�(+��'�\s�F�%0Q�Ǆ &(9�E
�������G��Mk�g�S�? ����Hܼ��1�S�X���"BN�	����DT�G�PY8���"|�F�%y9!�d5H*ب3p�7K���C�E���8�牊v�
�am�?�h��j�#^��B�I^k@��v��{}��s�U J���Izy"�'M~\rW&�DX������/|����O� *�+I(�(O��O>yP��l&T�"iR�b���(��U�<��dE�����%�Y�PD�pJ2�h�<A�%��z����l�#i ��D��$��x�M�P����W�BlX��D��0>�J>yEe&\��r�Aڰg+�Q���^�'^ўh���ԟ�2s�ɡ@{�upgؚJ�=k	-�	�G�qO��K~ZPf[�@ƹ��ϟ�>��)ef�Z�<��(��\�@R$^
�.�KV�U����?AC�W2v��,�" K�^I[�Jg�<)Vƚ/=�qs��dp��h�Θe�'Kў�'7Pց��$�Os�p��˓�o�TF}��'Ǹ'��)b���g�OZ�(���ar�<�=�����,s������JzCX	�Z�E���˴&-D��W�T�b�n�� \�#D����J'��|���O\V�&�1<@zS�j/��'w�12��Z�g�ണ�`���p�)R�r�փm����ML8-S���@�:�~���'?�>7mҞ4Wf�p&`I]O>]�([F��re0�O�؊weݮQ�ؕ`b�+	�&�q�"OPD�0�+2�|�Y��T�r�(%�w�	hx��ǌ��:�(���j�2�.�0��,D�<	tKǰt��زc�\�!�=�"Ml�ܗ'�ў�&�X�B H�r�v�{$ #6���E�>q���V��<��o)���a�DI�	1g�4 k�$Q�n=!� ����s@!���ʃ� &!���$i� z��Qb ��T! �B㉄F�T�����#���ꎓ�2���/���$l��PP�Y�l2�eӫ��~E��?A�BI��eQf�7�Vܸ#�g�	7��8�r���&��Ѝ���P���f-�;�y��̺<�
PY�F\�xi���/�
�0=��OQ6��!�2B�����K��yȓNf�1�5��44 �����L��O��=�O ������7��#B	�#���ʋ�D@�M���tn������ށy
�scWv3����?�ɴ>p����L<ْ	2!�Pm��3[�Q8�G	Q�<q��OpL� &//��<��K�L��hO1�t�u�Q=O|`UHb+W�
�8�"OLq{�,*M��*�'E�BX�A<�S�t���)��d�B߭Ŝ����2��T�kqO.�}��+X:	��hV�;�����(�ۓ 3�O�0أ���G]�v��6`��	�"O��k���|�H�����i�L�pG��[x�8Z� 7z�b��g���S�%�A�/D���a�E�����G�"}�ah�m��'�{��#E}����;?alu�BmM��y�~E��	�@��'���H�a]�TX"0v��)N���'�����ŭ-��Ǝ������'�*!�"b�J(��� N�_*,��x�oN�Plz��gl�A�������0>�M>���1�XP �T������jCv��@!g��O��yt.�F4Ҁ�'Bސw�&�9��Ĕ>�'�D�&?�K�LH2F�8���e���1D�pD��>eؐH���=֎�h�,LO���Tk�#N�zӄf���rw�'D���A�/,�cWǔ/le���FK$�hO���..����oR�HU��S� ��6UL�=9 OT�W1O�Px��O��rpjʃN�ZȀ�"Ę]�:Ap�{jq��� 6�W"t;�d"� G9�,B�"O�`�\)FG��KG�;�Ԝ:"O��#%�M� �*`��x>��C"O��͉�;7�x��/nl(rP"O�dA%L�-.t=�$!�|Wv	Ö�O�l�V�)ڧl�U�'a�, �mܗ4	r,��x���8����/���+��8�ȓZ �d���b��=��	�d���\W�u	C4i�J5vCR;�\��Lž�Q��1Y�ͱ��5bDl���xD��c�7c�+�㜪�B!�OD���'��� ���Hn�qz�,T�F��� �'9��A!b >:����	S��	�'���Q!�k̪����;C�
Ik	�'�<I)�˚�FX�UY�`,N��� 	�'I �vFҨ~xŁ�C5�H���Xm���	"b�A�U�=��A�꛱y B�03a�x��(B�6�������I�C��4d��@�NӴ	��SGA��	y�C�V�^�v�%6����0��C�-+�8��ʄ(U� ('���D�|C䉵`�)b�	U�iXtK).�d�>�OC]�O�2�q _	���T�H������'��%SQ|7ҡ���8!%!��'�h%���6��Sd�ͷ��= �'À\8P��ok D�$��8 ���	�'~ͻeJ�_���#B98Vؐ�
�')~��P)˳I�^V�j^ �ʶ�������!�S�O �l�W��\�pF�?8ˎ�z�'�
URS�\�sxT��aղx�r��'�nAkd��+�4���%Ȏi?�]��'d��� ̕
	��b�ݘL���ʓP.���Hӹ\�~�`iF�������&���"�Ll`�i��i;V�
�B�������X��F���(O��I>�#�>�,�_��ic��W�<QeMê�ܜq'�J k������P�<���	0K6�0��LR�X��b����xr�LiX�8�K��6?��(T���0>�H>�aF�*3jЊ����!Ĳ�1���D�������😩�l���{���B#,��=}�?OX�y�l���fj�,q��ѝx�^9���"��@��'�$�S���y(а�΂�9��G��hh�{� T��Z\�O\<h��P�ȓF!(����0-ʼ��6E���Ex��)a$�UO\�z�����b�����hOF��*�I�f�.�N+
��$ǒ(|�=Zꁍu:Pc��ʄa:q��'�^� mϟg�X�#��F�B�k	�'���X�fiv��"$���}��'�a7b1(l����(��
�'b�� D��?���cQf�w�H���)��<aU&�V���2	A��]c?y �h��h�����S}��a.�ldp"OH�V?N��S�� �J���"O��h��ۡC�����H�S��T��"O�X(�\�x]6=�H��	���"O��uFL39��f=���� "O���.αo�BT���J�TuL��W�>Q%,Lj������QF��Y4�	oղ�h:D��� �2b�� 1��B�?4��;D��J2B�2O��PE�7{�|�j7D�4�v	<}���I`d2O�d��7D�
B �Cr69�E���q.,��k5�OX ���'}dT)R�@�\T� y�Ad	4	{�'������"5n���*�*T�$K��� �����N�J��1���w@f<� "Ol�R���V2\x҇��!�;�"O*�{��S�<�Dݛ �O�d6R@zf�	B���)�G�a��Ȣ0�`�cB�\�Q����'扃����S9�n}��eJ�/�4�؀�]�@�1OvQؐ������
7�A%J�`���C!��30�؅ȓW��E���G�H� ]�ӊ�{���<���IB%4`�
W�S2$���lc!��3�ؘuFܿM��My�T7�ʣ=�O��O�5y�R	GŪܓ"�Q�"n����O��ѡ�c��?�D.��@�(Q��#l��iR�:_䠸��KAh]k"ՊW�dʄB��B;����!��1�S mA�t�Aƅ�P�Fx��'�@H�҇ n�0AH�d�䰪�'͢IjƄ�>��A���Uat��'e�	z���{@�P=9�!�Ǌ�0�B}��B���شSV��<��4 ���H>A'i74�2�g�#/p�� �k�<YE`�?��� 6���g�ڬ�c�V�<I�K��mrv�Cߨ�4��/G"s���z w삵6 ��7�e�a|�|"Ƅ4P���&�еf{�C�0?90�T��?	�.�6���(�ȉ8Riy���˟4a�q�OG�Y"��T�Gz���W	K_X��+�'�R��k�.p4��'�PZ��P�
ӓ��'���٦��i��di�&�c��R�'�D�e��)<r���U�=Zx�����$*�S���CCP��Q�T2A��e(��O�����Jr��D�؅a�r��X?�� ��X7qm1O�D ��=���K�@k�F��2\;���bs8Ն�&����׫�)��JQ@���<э���M����jӉ �L���d�d�!�9����@k$j�p�ACN J�h�=�O��O�����G��x2��X�.R8��g�O|�S1���d�OF6=���Z(l~���&�$�fS���Z��|��`�OR)?.��O	:�(h��w���ƫ�M$\i:� F�PFx��'��%a�G�i#��z�(w���q�'Kѹ��B-L�����v�>\�'��h�����H�}�����h降	����o�? �F��<qǊW2 � U%� g��iT=�6AѶei�Ua��'D���f�<\g�@eĊ�|�p�`%D���D@~�~�`i�8o��B�F D������'l�6l�5oǊT2ud?D���T�ݚ?<�L�vEڵMq�ѻ��;�O�a�'~ة�a�=��l;�`$,ј�'0^�hÅ3]G���g��Y��I �'�0�Zs��%,vD�� �e��5k
�'�)c�'H�X��x�g+N/X�9��'Q:�c`I���RD.��V#�D��'�<�2�N�f��qJ�-�;A �[��$���>9����4�H��ڡ
��.D�P���ō4�Z��aN� �еS��.D�(�6��>UJ8��	F�O����0J!D�P�։e�l)�.������g D�s��]7:T�P�L*FV-B�
?D�<�E��5����f8^A���O`PJ/(�9�""|�ɊJD�4Rf��9X��d1���hh��!o��p"u�>��yD�ͳVD�à�1D��IC�ϫ6�8��@,ּEt^e�..��<��Нn����&D�(D�[n�<�!4sO>0��iO�P:��@&��<!-O��=�L>���5���.�>�u
�gC?	")F- �GyBp�I$�I��M�Y��m�$ӂL�B��.S!#P�X����S&j��F�4B�)� <`ҥߴD����(6^�u	%�*4��f[�}2��Q� �1*^��D*�OēOvM�C���o�(����e�6�����b�'� 0)E�'dv��aV*u������,O4	zJ�8��ڗt�\b�0��<�i�,v�,$�d�Ƨe�t{��R��!�$�5����I�4.%��#U
��az����+��� /����сH�>m�!�DD]���g�$Vf�H�=8� D{ʟL��A�:l�M�'�5v�����%������yr�Ȫ��T��0'&~� bÿz��ᩔd��'T��9��_�g�	�M?.�0� *��GJ�}��B�I�=�Y�*�!x:� bfL��b�hE{��Ł�!�la�+Ƶ|�jٙ���yRhR�øXaHZ��F<K��ҋ�ў�'��'R�D�%�(�Y!aZ�w{�e�p��p���O��$�PR�Ŋ���O2�d�O��1�r�bA��"1$lXT������0l$ш!`��O� ��T��J��K?O��)W"&zr�@�ЩdEM.U����+��Ly�c50X36��x��m y*��	��vũ���EL�D4?�cߟ�S�4�>q��!��Y����&e`ìCJ�<��Q��P8"�؟z(Jx� ���<��']p�����O�R��>����(uʹ�ĉ��flֆ�X� ���/��\c& ��y��OV�L�@���	Bq�x�$��ذ:lܫt�JLQ%@�' (�SL�rx�(���\���H�����m�Ţ�&,���v�@�dqb}Y�Iox����̾���&jRR�`��Cҵc|����OD�=	�}�/�"AʣN��A��0>�L>IAE��N�f!���R�`|�)s֤�ZܓA+�Qb��������lz>1l>r��S#��gC��H�t�����$@���	�|�Ň+�p'NI&9��$�
~F��ԲeV��8����ay�4Q�p|�"Ǥd�ɗ;b��.,s��UQ��B;�����X���'�I\���O�,t�歙�m�b;��T��Ɏd-�Qz�%�E�x�B����B�i�L�YK��a�ɪ�ᐅGڦ+��ߟ��';�=�P�����'��Om�Vn��f�f�jGˌ�r�x��S/�+��d�O�P\D�P�];��1b�O�`�d�ҭ�"��RL�n���jd������du�6Έ8R��˦�Q�2�$�x���0���b ��S;v"�'��>�nZ-G�^Ȩ�B� lG�A��[��B�I�,i������I�����a� JN:��ĄK�'�ΡJ�Nԫs�p$j�1O965Z�'\�`ȁ�d���O�@�&F�1s��/5D4ѕ"O�`.ǹh��	�ǯM-2�@�`c"O�*��P3n[�l��ij�I|x��(1	�
:��8j���+5�h1�j:D�<JB�=���Q4�V�P�V)Se�8�Ii���O�e9#��U�|�����0C�4���O�6-XU71O��ݱ`QT�$���g+7
P���R璶w}�+�):D����+�	1�4��f�?C 	85-D��{�G#�xh��-FڀI�g�}h<y�-~��r�H]L� �[w�m��&� ��N�s��(�J��=2|e�8��hO��#���O��)7��4�fe*��ʠ��ib�>QgoM�Ak>a�<A�kS�Ӻ'�ub����U��P��|> C䉽fD<�4����t�f�Z/�����+�	�]U|�C@3;!da(��M52��B�	�@���ytJſE�0a�A��p�"<����?�Z!���Kb`��咏dp܍C�Gj�'��u�Q�D��yw�Ս9Vb)B�C�E�3��=�1O|����/����B�Li0ƌ�u������R�e�ȓg�<��*�`o.L�t뀉&x�<ɍ��)I�����I6Y<$�� W&�!�$ښ]�Q�$�2p4��B%H+-��=�O\�O�eQ�IM�0�xԘ'�J:]U��A7O���$�7� 4  �   H   Ĵ���	��ZZ�GbO8;�TY�P�H��R�
O�ظ2a$��X- �F�i8�6��,V��	�%�X9��2�
QY,�nZ�M#�i�V��%BM)K�A��r@��i����8�OP��M���O�O�q޴~�͛���4?�\y@�+Ш�'g���`��E�+O~��U/͙�� *O���tLz=���G�/3������?%���e Q2�?!"�'n��`צ���tγ<�6�ְ\i:�)�枦 3����P'V��FiK�#g�㞸�D�7k���+YJb���nW|�� �r�E�B	�'	��Fxr �m�	�)C�	���l����iN���I� T�L���	�IX�T� #"�����	:a��)x��dC��Ozl��O������(3��b�I6[��̓a�>�7%7�X� �D�E�8мy�Γ��+�al�v�0��d͎�O��!�2+BV�(���Q�đsN��)_�O<�k��d�'���ˋ6���փ�� ���AA��x&�0q��6���""Q��P�Z����.~40Ѝ�d���O�+�wł��e�_�݌�����Z���<9�J*�iǦO$Y�����r�kH��5�8�9D�Z`?	U.(�4O2����'�����%�p+��J�.�����ŞcB��Γ&���#̈�1ߛf�>�B"Kܺ�t�'������T1�F�@�:++��*O���ch� y�1OĀ@� ?��J0R���>�k���8aL+V�HA'�I,)�@"�(�ę�iB�F	sB�#D�8���   �
��W%.�@щ�"O�q���ٸ*�b�7IA9�M��"O�b��S6��)E�oU,��"O⤩cW�>r��33���:U��q1"O$��^���'���!���`"O�h;%��	Zx1����R2ꀓ�"Ov�)�CW3~�X�פix��"O��+WL�jpf �'`V!ش"O��[%I"Z,z�r��]'*~��[�"O^(js�A�Waƹj�K�5w_@�90"O��ҁoǑ`Y�E��QL^\�"Ov��C�ΡQcl��A蚔:IXȺV"O������ �^�a�fY�~4T9f"O��G+�/j^,Y�S��P�r�"O���Lҕv:ݸ�\��j��$"O~lR�K��^��:@ 62:��Q"O��I鎵 ������:3H`s"Ob8A3�� [���U`� ���P�"O����R��4���n�)    >    :IZ@-�nkZ��&C�'ll\�0�Oz+��AI��e���X�'M�X   ���:&�4����6�ƨk2   c  �  w    k#   �pA���d�Zv)C�'ll\�0BLz+��AI�o�'�|)��>9ā I22 )��_�nhr���e���F8��>�!@��-��is𨗣=.��!`BW�v����.��>�1)ЖDuV�v�ɧ.�����ߣ-����&��	�H�>q�.hM�4� �L-���TZ�<�R�M#T�L�(%����h��W�����'��O��e�O�
-���!iW�u�6 B�4��4�
�'����.�/Z�� ��\.<N��'�0����=�R���J�'*��"�'e&��%�e�4a��������'*���0��;t���A��b �;
�'T	���29|�G<%� ����N��>��._Y1�!����59}|�B�'D�hq��G�l�"l��n�D C��!D�c�
�e�xx�"C�a`�� D�D(�FO}n#�@U�E��r�2D� +'�z|�M)ÎF,b<X\�F1D�XB���.��R2��J�\;�`����֊+�S�O�f��7
�9b\�I�+���r�'5&�8�˝7f*`P�J��V���'�vL��GF�U����>I.�Es�'\�Ń��3 �t��18��]R�'z�o5"��	6荹Hk��ض"O�	�)�..��+&H �2�8ڦ��6Y�Z�Iq��s� �!X��%�DM߽5U�9��Ea`T̃��Ox����הw��@i�l�#0ss�^`ߜ�xV
�Ix��phTB����ƆƖ��b+^�����O��D�O���?a�}2���6$[��V6}�A���y��9�� �pЬ���:a���'��6��OR�@[���������|S`j� T/f��:�"OF���]
���e��Q�H-�t"Oh`���̇{9�y�vʀn��h�"O�9�'�L� $Z���)�X�$�"O������\�����#��5r�"O�p鱌	,�d�E'��$�[V�䇈
3�=o�V�O�ZM�"�MJ��u0c�Yb[p��L<� �+����O��V�U�"�Z�J[RL����K�E�I��Z��?�~�E�A�CW����sd<�k��C�I#3���$�O��������$�82\$�J�Z�y�xp ���O"�򤗖~z���X	� ��I(D��m��	!�(O(���o��p�~UPCjP6f�(�SLw�`�IKy¡�Z���dS2=���C#� Bd�d��$z`�O�e�t�'dd���K���*T#W�S<Rq��}b��<�C/�5��|�c�����'��܂#���0f��L<Y���aZ5�1��5*�"��SA\�<!akֻ{��U�UɁU	�Hr���T�DM|�����xIٟ�����Jū+*�(oP�"���Au-������ʟx�ITy��'&��'@bt�B�S�dIa��MJED�k"�AE<ի��f��ؚ��J	� 	���"p<���´|P=��"A	PS����?p騒�vQ��f6YK�!�O���WU������k�@[�����¶Ul!�`�����E}Bj��h�
�q�T�I@mؙKbZLc����O�5oٟ�'��|�s�y����hӨlb�Ĥ{JD `�ǒM��LԄ
ߟ�'.��'���&|R)��EW���I%�I�rN�&y˔(f/�%,����խz�\�a�ڄ|/�ɉD�4i����%�D�r쒧_݈��dw-��x��qo�⦩�a�U.>*��8�.^�b�����m����D�O���?�
Ӎ��F�2EXh�����%�x�А{��6�(a��1q�Pv��<��ǭ�d *���?�(�ʰo�Ӧ-a�H�Q�c��˅gvb��TВ�?��.
f�Q������Y��*��_/h��4	!�S�^:��v !�D��z�!foeŦp�V��O�O]^	0t�°'�L�zd�����|H<��ş����ħ�ħ?و<1O��q��!B,� K�B5�=y����<�5(ϿZ��D�K� �<��`����E~Cn��YnZ{��B �Q�S��B��\[�� ��I#]����?��g�S�? j �v%T�G���F� P�R%	�"O %���J���(	�d_$��u�"Ox,�@ɷ/��A���SV�`��"O��S�I݂Qjd��VU��@"O�8pc�\:�Y��@�~5���"O������9)�܅s�BK*�����>��Zi��l B�ةJwv����XJ�:��&<D���E#ϙ:�� ���_3N-�6m,D���Wj��3����AC��l;@�.D����L�G�$H�(��2G�IR6�.D���
�$<���2V]3tc-�O� ���'�����6 >�Uh�;�f,j�'��e�5��y�n��$��4�T���'��hyt��>UO�0-E�=_x8�'5��9�C�3&�BA9��;5�޸�
�'n���'�MW�\� �
�~�vY��'ƕ U�@6'��Z`�Ƌ}͢�����-��>%�`�P2�NdAD�4ȅ��*.D�$�+R�!�EK�o\!o���H�8D���D�T�0Ą���C�2y��A�.4D�4x�	�m�h��îؓ?Ԗ�I�+3D� �en�<R/�I���W�|��-ಆ2D����L�;>j�%�s/��etdq:$k���4�>�S�O��H�e�mv�h�ʚ�`+�'�f�L~��1�[�P|�a��'�x��F�ҔH����A�S8 LF	�
�'[���L�J��a!Fv�X��	�'@��:��˺VD�R--n����	�'��!��O"x����{��8J�+�F&|O�A���˺��UKR�Z��2q3Q"O��l %v����Oмf? ���"O���@D�!z:��N�9Q:d�*c"OvHEMN�Y�*���I	%`��""O hqVLBA��Tke��j0�̈��'�\	��:�h���%��u'��	5g3:�؅�ȓ�.���aϻ6��ęaᇬ"��ȓ32�!���d�\8��I+����ȓAf����h��hk�)K/Y�P��Fb�"�!�D�f�a�`�U��Ѕ�8���Uȅi^=��O_�}hJ$G}2���h�.�8�F�8��2�	Vp "I�'"OZ젵�^%cZd�
q��;P��@W"O $�4�?Q�4�H����m�L�8w"O�a3�A*�b�c�P1iӺ�U"O<8`��73r��	�- ��	�"O�U��G�B*:p��e�!\�L�U�O�&�)ڧu�,��[wnձ��^�"`��M�&\AV�Β�2�����!a��Ѕ�"��A���>��������F��z���G1G"H��C�	MU$-��7x��2D+)0'����2+�ՇȓR������P]��ВH�;2jj�ODuZV�'ņ���$[�!�*��|�,,��'��mꥮE~�-�2�\$-��'��jBDH�lit�B
��!G��p
�'Ű��e�I8O��a!�G 9�"� 	�'
��:��FBY4�9C`D�Fe�Q���+���8:��`K���x��%��$}��C�	19��ek1R<2��S�W>,��C�I&&~���ȇ�`+hD"��ց&�C�	�T�	�蟖F�(�!G��+�:B�	=d��� �F�	��H!1�M /��B�	6��T���o�L'
�8⸢>�䃓J�O��X�Q�]�B�i� -�/
hQ�	��� �AQ���V�f��� ��(j=(�"Oε8#Ɉ@��\�� �&���C�"O�����|�ơ����
F�̪t"OHd��۞�q'���)r��"OZ���&��Z�p1i����v�
��7�Oz(�s�)ڧg�p�#z�T`@W
_  �ȓ%Tv���	
N�h X�[�l�$�ȓ5 ��q��l���;�ڜ2�R���jod`1CQ�O9���Nz�@�ȓ2"I��q��I˱j�dV@���4&�}Q�H�d����
R��O�b��'l(�F7����dT"�`�	�':i�Q���H��b�m��l�4	�'��3��Υ4�=@w�Vx�f�A�'w�=с�W�;�J`�0i�����'���2 �.�d`�Dț�c�Y������IY�9Ss(Y�FTZ��1 :��?�lX�򡘎�l�d�I�2!�n|���ˋ%1�����FF�%.!�3KM	m٭�J��&ψ/!�܎�(����YJ�6��e��k!�$�6}��-g	��xPt��e
VQ��(�' ڧr"�"� �� �h���Β&.�t�ȓY��1��D�~hA�r, '(��ȓ4 zbʃ t��D�C�F?l��>h�����%!��9J�
�*����T��	S���b�QA"ӭ35n���"��y�0_,)sg��Q@���!�V}Fx��	�1|e̽�u�ݝ5>��Y ː<S!򤐸n�����u,�� ǬT��!��l��HC�@<Z�������!�dG�-���L�6)��D'?�!�D�&��E�բ�K�(  ���]�!�DFg�(<�@I�j>�YBS�J���t+����ɜK��±GJ*�t�-	)ԄB��S��Cړ�dy�n��T�VB��8b�]I�-Hn�|(� ,�1f8C�I�J� 1�M�D�p6��i@�B��<^���F�Y�;�>E�4E�F��dXn�.ɫu�r��v��+C�Ȱ���yR� 3�Nq#�3$��|��gB��yb��Uj&�30i�#��Hz2�ޒ�y�H ��Pa�.	@���y��.�����`�A�Ý�y�l=#�P��p��� ��"a�C��O�-ȅ�&~��� Y6bcu��? �`C�	�w��A�
�<�&-��KP��JC�I�+3�d��iA�$ 6 z��ΰ��C�	�pV�`�
C,
p��և�zȘB�lY��F/�Vx4�H�́�&�jB��ȍ�Bo �$`���?�,�����#<E���{O
Q�#�z�>Q�3�P��y��n�uR�N�:vPB4�"�_��yR ϑ�V�r�@�}�Lr��I
�y��	*Ӭ�A/|���@��̈�y��[�z�@C�֮d��ȦBL&�yB���L%+UI\,,E:%	��:��I'�t��D�,Z�PzDm[�B �H�c�:4!�h7.�PGL�6(4iDd=�ȓ2�=i��Y���CɊL	H��ȓ>P>08��E2&�h�2m�̖T��W3d:��Y<�XyREcۯa��P���P������}�x��c�=6�#VIEX!�O�\ p�fB�Y)>l�4j��E�!�� 숫�
M�Iq������m�4��"OD�bD&/>����y�L��"O� �'�NJW\���*��0�0P�"O29[fJ�|B%�A�H�x���#�IYj�}�� DZ�y�Fg̑|G2I���u�<��c�־�
w.E�
b���C�q�<qW��`(tp�ǇO{�9�t	�f�<� 藐M\�D����Ŋ�e+Nf�<yq�ܚu�p1�A1L�r�B|�<QA�O�IY���B�:IS�ѱE.���1��;�S�O�b}��mT�k
2�
��Μoⰽ�'/~H K�$42+��Ő�(�C	�'����R��7��b�%�����h�'�DCf(��5P��$�7 8��'T����{�MJ�
E��)
�'b����'�]�)���|����I��ѥ�:|OJ��hG��$ܪ4��`R�"O�l���� ��1�`�(�C!"O�@i�F	s1�YkS.� M�,�T"O��@�-�`�tEil��jx��&"OQw�Ŧ>4pĈQ�eٚ "�'�vu����M�#�_�z��m	E�Z�'|T�ȓ(P@�׎Be�I�ҬUh⑆ȓM� -��?\	򃓁-O��ȓ�r���U$�A��.�K�<	��7�uN�4x��g�WS�<��ʌ'G�@0#LQ�F�� �!-�P�'P2����)���E�d��$dMz�"�(OA!�϶i�z,2���1&*f�A��W.^/!�dƢ=�X���K��|�@@	#'!�DZ�H� m2���D�a	2�ݩ34!��^~c���Iʩs�VT��-	u!�$>T���i ��z����I�t ����'���} YW�`e��B"��}��I�<��[�-��\��&�7#�6 �V�I~�<)�-�Y8�E �6x��	���z�<9W$9e ��8��5X�dm�0o�o�<iB�ݒv7Tp��J˪?}�����n�<R�»��$��jٕH �]�1Ɨb�d
Tn�{R��+M�Hs�RCJ����A��y��Q��h�C��X M>x�HE��y�a�l���"�["p�T����y���ro��2�n��i+h2#$��y�+�
y�$��7��;R����� �p?Q��NПk!�÷ʲ!�r�ӱB��X"�/D���3/�I�N!8�k�3Jޤj-D��C����"�\�;��dGxu��-+D���2OE�GO�A�r�N_�|�*��.D��SS�	T��-�b��=X>̒��!D��v�H#B�m��ғ?rh�*A� �r�E�4�G6� i�N9�^ �됒�y�MɊb����a�	,6�T�� �ykT�t��b�啒US��ic���yr��8O�
����F�a)�|pq�\
�yRcҍd�횟'�4h��F��y�]�x�Dy-R8&ʽQ�aH��~���O�>U:��H�^{ju���E?Z�R���$D���F��Ƶ��K�C�:��N!D�|	�bN�:Hr��S� �f.��8��$D����Ɍ�Ur�lPB-J@?����#D���o�p�p �L�iPT�F D� Rj�)L���Aɩ	R���6*=}�\-��=���*V���C$�%O�X�00�]o�<i�8�P%P��\�I#i�co�n�<� �:#��C�=��q�$L�2"O0��CI�/Q�����D���k�"O�,��b¶P���C�.��jS�'R$����%�
��r�=3��S6|�ȓlN���I5�j
M��E��^��Q�W&|���cQi�̅ʓ#�L�j�-B�zH�"e�-��B�ɛ,Ƒ�0 E�91*h�B��!r��s� �"mo!k6��8�v�>�@��F�O�f-�O�D!"�H��U.�t�z	�'� jrhƨ�L8Ŭ�
b����'��D!�B+dPc�R�>���'�~�S�N=�j���݈z���'��ei����ؗϞ�p-r�I�'��ɒ	�9� x�BW�5�]�#��l}2�'��/�s����?�����MB\I5��B�[�\�)���'��d�R$��Lb.9����W�g�-l� ���W�M�l���"8TY���	;K��G�'#��YA�8�3�d�/*P4:��Z/=��p2��_�4��o~dL��?�'�?��}b�d�6��V��	D$@�5�P��y����լx3��O�7���*՗��	 �HO�i�O��j�
fk
�N m:qɋ:G���6�%�yr��p=��21�z�*lXZ���߾!��Y�
�d��E�E�X���<��U�]<"l�1�ъ(L��"��+�ѣ&%�/3�9C�	���<��1R4��T"x�LQ��h�����F{��$��jV �2��]E2�x9mI�����x�6�yPL�%8�����A-��'9�6��OHʓ��a�QU?�mZ�h�a��ł�8fV��$�R*Pt������Ol�$r>9ȣC�"�ґ�E�y��X�{wظ�F��� ڀ�p���<���/���C�3@P�^}�$h�w�@�?p��ә)ayR��T�D�O��B���hx G��l�^�)��)lO����F�hp���h-�P8V
Ot��I��x�⍃9O>su+ĕd.���<��h�?�?ͧ�?II~�ڴ-���E�G�e	5���!��ڂ�'��\TӲ�ڏ'<>Y�g�>�O ��b�RXBP�1F�������T=�O,� �� �Oƶ�Q�R�O����VxA�����4�I<ɲ��؟��	y�OЛ��U�,$��s&�J����Q��y��[S� Ċa!V��Rĳ�	��p<��割jD:�B@ /^�v�B��Xo���}v���?I�g�+� �7��?	����)ߺV-Lهȓ&]�y֫�eMJ9bVk ��bL�� ݸHE�Y�B�Ƞ��a+!�lD�ȓ9��L����7�}� �T�C:`���E���n¯Bc�YS���|�b���AY8ӣ'O4g=*E����A�8��O��qW�'�(�x��**������!M����'��@���-��(V쀮sy�� �'�\���b�[S��Y�Ҥgm,4	�'�r�vi�hVf�2��jE ���'���"�g��<�ޕ���Ƃ[(n9�$�>��	s1f\�`��	XjK�ԷB��B�	?yv��T8b�&u�c�Ϳx��B䉔$3|��R��)'5�RwML�n�C�ɖmm�����J%�l�?:VC�I&~�ui���R��Xd��5\�xC�ɣ8��{$�WOÀ�vϟ�_.��>q�.�A�O�b���'��Spxt
q��'#kP)R�'K��V��h��b��"f%j��':]�fn� ��u���fӊ�C�'dr�%+M�6:�X��i�1��'�;Qm�	R�Y���:	�9h�'E�ɡ�˹{��QbNY�`)�
�'R�-�� ��   X   Ĵ���	��Z[F�ƈ0Z��SeB}"�ײK*<ac�ʄ��iZ(b� @x�&`�,�mZ�_ty���W5hR|H���.tc����4-\��z�l]��	7'��$����>1eV���DT<~[�����ab�'.�	,a����ճid��!�BP̛D�5G,�b�O �ю+�M�4[�8�����t|��SU��Z��ݕ<�bI���"�V]{Q�݌(Jp���/hJ�L�O������uwğVy�aδ6��h����&wd�JWgya�˖�>پ����`~�J }L�l�&Ǹ'�Ll�H�$����yǚ�JC�C�BiV@'�8I��'��'�&H��oљY�H#��<}���'aFxbf ]�'-����d���R��U-RԄ���&�O3h#<�䉹>�FLD�W�Pl��-��|�~�i�O�`�dD��O����{r�
u���S0M��F���M�n,T�*"<A��O���Q���-��|���V�p�`q�>Y��#�`K��~sD}�bh¢|[L��倞�G���'t�Fx�A��:B�I%��|q�jETG�ѧ�;�N��#<Q���O���ʈ�>�#cjPY��(9��O��O��N<�'���ʀ�sO�= �������Q?P�3~ 4O��@�F��9��	�@E6PKfG��F��p�+ra��e��9U��	�V�>	0'��,"��	P���@��l�"�Ë�	J�Nʓ���En�|��$ԉ��3�DϿ_Y(THS����	X�$&���:���������ѥ��D\�(yV��	9XB䉘u7��  ���"O�T���I>/��S��A���"O� �m�4�h8x�B\�l�ʌ�""O�I���_,|tI�D��6y�Ha�C"O����xZ�$C�Oјm���[�"ON�8��9F[P�{�o���T�%"O�	�`��$M�@�s�O�]�fe��"O !���K�X����!-��"Ol$�Fh܉r�S�/%(�@�"O�I�D���M�b�Ey��XY�"O*��Ջ�)Lǀ�j�ȎK���Q�"On�%E�_gP����	k�b�
D"O$���W7tA��F΢/�$�Jg"O�DE��'�~�!� ��4Q�F"OT p�dC�%fmj�������V"O��c���_q^)�1J�Q��	7"O�)s�B~��YB�f�'_�� "O�<�gƗ!br�Qץ��Q<<*�"O�E���9-t   >    :IZ@-�nkZ��&C�'ll\�0�Oz+��AI��e���X�'M�X   ��"OBx�DMFU�{���   R   Ĵ���	��ZDZFI�>C��SeB}"�ײK*<ac�ʄ��iZ(b� @x�a�,�mZ�|8@� �>X��cYD�V5��4j[�FGo�F���	#'�ݻχ_|v�
�Q�ۤ��^<V"��
-�V�� p0�iJ�r�!ɌC㢤��*C#t4���O��� ��9�M�G^��QjB�2$
gR��Z���8ˈL�����tt��v�V�8�H�ÈH|^D�OJ����G��ugĚSy�E�&t�� O��v��g�Ta���>C�a0�&.?�v[ }y6�\ܓy��ɾ����1M��m��M)"�N�AO0Lэ����mr�0	��E* ���Hp�ʕw�����#<��*@�^�2.:�6u9�׮A� �I����ʇ_�K�dL�*>�5��.�7���t2}� �I�'�X�=�e(Ֆ�"��'Έ_m��F#�ݦY��I+��ɓ��1Kb�<��c
�G)<B����[��b�����ɥ2��	�R%8 ��,�hiat OT���)
N#<�$�>��^���	pD]�~�F-�$�X"O���u�|C���p�'�*�Jg�U#|�p����+��UQ�yB�[]�'���$�����$^]��d
�h�Z����" �	�[��'V����>X:H�ǣ/c�Y�qN��"�N�cj��2�	�g���Q`k��M{K��;'%w����e��$Rwb_�'���p��pWTe�'ȍ8!�×�')P�x&\n�I�V�D�D�����Y��� �"<��;�5Ἤ��Ӹ8;�P���+Q\@Մ�IT�  @�?��
�ąR�"O���S�߮|��,���53�-�"Ot��%F��q���R���lbó"O&���m4r1�m)uȒ�*M
b"O��"b�P4|����$9�iu"O�M�� YQ�)хFX�Ov	�"O ,K�o��6�0��ЪDl� @� "O��Rq$�<��eIL�j=�$ �"ON�+��pN�-�ŇI/��5�e"O�ÒJ�+'���D��0z`�"O�����G�ޑK`iA�^_�	h!"Oh1"ǌM�
��y�EBL@b�YQ"O�u�"B��3�6���f�O4����"O*9�cõ(PZ�Sϑ("�i�$"OR`�r�M�:d��M�	��qc2"O��`M��;���xūC h��yF"O��0-I�vG� �qJԮD�=���t�O�t�aU�e�ꄰ��X�}8��C�'��S   >    :IZ@-�nkZ��&C�'ll\�0�Oz+��AI��e���X�'M�X   ���*^4��'�Vds�d��6I"�$O�S�����'���R*]�}������ժ2��ԇȓ5K���c�cTv�0�B*8�,}��5�Q	ы��$n���,&<]����$�&�AB�Ǐu��c���aHM��L�z���Rk��BA.WW�j���
/x`h�m�M� �A��G%i��(�ȓZ�����K��tY�{ԄѣPɆȓC�5Q蔜���F�I��"���h�PǄ`C�r�,�^���ȓa��-Å�
>%bq%aJ0\�����}�$o���0R�Ƅ�W0�%��-�N������������Q��X��/%�@P@�ÅG�\�	��0K�I�ȓxX��eٿ-�~�C�,U'"2�ń�vB��f�C�u)�zs�:Z��S�? �!�U�B0.Ԏ%���":�qa�"O�E�U*��%�J4@���<>t��"OL��łS�}� ��n��xt"O�H��̋�M�2`8 "y�6l�6"Od�sr��eil�P�Ob�l��"O23��+��u���](�V�8v"O��k$�ǵ ���ke(�z� ���"O���q��Q��JC؁>�Ե"O<!cB�߶#��p�&��Ljμ��"O��I�铒��0ȗ
Z��[�"O�P1*	3�X\#W-�#����"O�ٶ��tf�e�ŗ6r���a�"O�	����5:��t�A$R�}p�r�"O�d��*�IE|��� Ib���`"O���BF�X��z2e�U@t)a"O���SZ�HDɩ��Z:(!���"OH�#Rj�?+�XT�ЁޘC��q0!"O�1@�d�1_���!��C�j�A3"O�T��'�%Ǭ�I� 5-�*y��"O�\!e��.eq��d�Q#��T��"O�aC� ab ԁ�ᐯV8e ""O�Hq��\�TĹ.�L��m""O~�[�f�n͔�;��6g���!"OJ�c���w~��Vn� 8���C4"O�g�W�4���Z3t�d@��"O�T���A�F*T����Z�}���3"OH�0Q-
w8l�$˅�Ze��"O��[S@��[:ܺC.y�	�"OԼ "��~`<F�3?���"O�Q�6N�*�T�[v�SD:���R"OV��G�V��w!��;4-��"OR�23@���f���"O�#
\/w�؈7`6/�|�¤"O�5�2"���1"�F1u�T�%"O�e)W��#b�0�3�./	� b1"O<9�P�Ξe"i����mx@3"O�X�f��|uPa[��<5rD��"O�e���%���s�ƻk�*�J4"O��V���H��1��I���r"O�-jѩعoS�x� B�ڊ��B"OxɰG¨cL����R�k/��0"O��� Jb��MHE*a"OL����H�,pL]����z0�ٴ"O�����j&�i��{ܬآ"O��#&����=��X�&�K�"O���bA�]s�m��3��"Oj�{ѫ�D9�)�AÎF#6݈�"Ol(���94)�Ɇ-�@�"O�)��5;��I@�bաk	bst"Oj��H�@��h���LW�=8�"O��X��]'?N�BA>];���"O����9V��=�uF
 ).@���"OJ�z�II���l�0�6&,�(6"O�I��L�*C.���É>F���$"O�������TJ��߫H1@��r"O�1��~�� �5!(s��$"O�x�a�R$ZѶ�H� ��f����"Of\RC�+i�8<�O���"O�Lq�N�@)�A d��	@Z\13"Ot���LK#]�p�a͋|9*!�"O$(w�/'b�[��O�$|IҒ"O��`aX�\F�(��*�~t�Q��"O%��$̔�3��F�n�p�¦"O�-�PnW�1=�<J�	Β!�&�a�"O� �q�r�� dJ8��%�Srb�)"O��DMϪ^�hС4g)uU�h�"O~���H9�B�&רT2��3"O���Rj��s҄���˵Yi�݋�"O<��P��0�2p����p��8�"Or�R��׭����i�,}Ӯ���"O����g�U��H,�B2"OR�z��E=[�b`��B�+�~}J"O��D3נ�C� ԁ3�TI��"O�uk#m�.:A�F�1J���q"O4tP�%ŧ"�����o��NP
`"O�qA��K>rPTX����N�R�"O�,ǡ���aծ[�\�c�"O8��C	e�8=�N����1"O6�!���N�.aS'M+r���"O�9��Ě�s�><sЏ�,pp(�"O�E����`x�͸gOƒjhJ|p�"O��#a�[F�$z�lO�_>e��"O�a��+j��a���ĖB�	s"OVdS��Nf]�5M�e.�U2 "O����M7�<�i��F��a��"Ov}�Ц�92��i�Ɂ�J����B"O&���aЈre��k�ʗz@��3�"O� ���Ԑ8�,Й!'�X��HA"O
9����.t�6�Bv�N$VQ��;�"OD�kt�O�v|qפ�-VK��A"O��෣N+B"��Q$�;b24 �"O���/V��9h'#�"�|0D"O�@S���[=�٢�B@gԹ�b"O�x �дJݮɹC�U�<�W"O1��!���,m(vg�5��2"O>4�J�L�X��v�]$f�P�bd"O
���fW�:��� Î��L�(\�$"Of�jr�^�N�j��M�%Z<�R"O%��*\4�\u���ti��7"O��7 �/E+l����%3@)�"O�"��*��5�2e� +G�|��"O(�� '!
�PZDIڬsL@��"O(9��h�_edġq�t�r�	�"O
����Y0dh-Y$�ʰ}��+B"O ��(Z^���ɉ$	h��7"O� �d=u���6�Q�>�z���"O,������`�&Y��T0K��]s�"O���#J�p`�������u"Orh%��x\`i��D�x��B�"O��w�α%*�,�r-1]�P͋B"O��ôjك$HD��J�aR7"O�&�[�ջD�.Tj�c"OF\�f�Ww~,i�C\� e4���'��U{D�I����V���,��i�'/lj��\�z@��"k-%��=��'���Pu ��b.�=�Q�;g��)�'�I��퉝v��Q�_�XO��'���+�gp�	�/ʗJ8N���'f�,�1拓?���"��)n���g"Oƍ�"N��w0�A!E�0�F|"�"O�P�R��%!�8�B�c
�<���a"O��@я�8kF�K3"Ϝ���"O~9 (@%"۠LB���K��e"O�zPρ�@-x�ke��A#�@B�"O��@��@ߎ0��lω����w"O�D�OT<'l\�b��	z��I�"OD�`솃W:�d���i�����"Or��5�U=z6����/J/�X�E"O� �tĪ{��'ON";V�z"O��P�:_݈��7�A�"O���uL�:*��Ⲯ� G��a#"Op����%� ����Bz�� c"O�X(։7|kT=���ݘ=�^��'"O�-ѡ/�!�X��a֤D6$E�&"OXk�f��5����I�E�"O�p���'S3��0��-8�xd"O���2��r~�b�@��\�,�D"O*�����JN������29�@%�"O��� ۪/�cc�G!F`SQ"O��"T*�.�n��aOE=8��T��"O�4a�ǈW�cBn��z�aK�"O��ia�<_��iz�ҭ�4m��"O$%� �	y`~Yv�A
Y�\�8�"O�K���<J�E�&�	�}��"O� �4\悑�&#P;�� �"O�HRa�J�c �yE�[�h���Q"ONm�rND�62p�'�c`�hG"O�0@��
�� �"L8gVa��"Ot����\$���O�|e���u"O~���ʛ7"tD4D�J_h9)"O�}HG��+�\t���=[d0)�"O�9�g$�o�����ȻaG�Ct"O���L4#�6%�'OG"��"O�x8+P�&q���I(�5A�"O��B�� zsb^M��y�"O�H�`B�(�f�x0`K�'U^r�"O`Qv����J�ƌ�%=:�5"O2���4[��t�m®jҒDأ"O�$ʦ�R�d��D�`��7;+樰D"O�h)2��t�4�/�.A'68�"O�t��m�.BX�N��'����"O2}'l�:L�"��Sm��H�ր�%"O�X��*̶vA� *n[:"B�"2"O�q�6瘗J
:�`۪S�,��"O��+W��(9��",�
z��Y�"OUH�O�@Ss+\�,Fn� �"O4ys��O��h�cZ�7I�H��"O�Q���ȅw�^ 	��Z�bJ���"O�"QW2pA��
f.Ν4 �h�"O�I ���0W�8�:Í7L �`"O�s3Ŝ*{�t���ƂKЀt2�"OvP�1���Y=
e�ae�d��YD"O@�)!�)y�aU��@H*�
5"O�h�5gP;I������S4%���"O��	w6A���r�/4Êh��"O�q('+>P6Z�R��>U�z��"O���&$r�jt�D�A���0�"O>��G(���ç�1Z�$��"Oa��J4�
tc�"m:�Rr"OB ����1ve�Q�A�(����"O�U�#'K�;�ɓ�F-���؂"O����N��Ȥk�/D�Q�*)�"O�q�u�D*@����MԜ~�K�"ONi��K@<YF��6�J�t�B9YQ"O����eB�R���wO�#8|�T"O�znߘ\Sh�@̾p!R̨s"O���5��0n�ȋ�Fi�P"OL�$�-r�6����T$UY@"O&|'�I'4m��7�ϐF�X�"O���cI5]�ڠ�!Է"��{Q"OX��
����S���<�L3�"O"8A67��ak�K=}�v�a"O� �]�FB
��8"���9u�\(�"O ���'ev�!�@E$_ڌ�&"OB��0E�d��(B �"C�>���"O�����I,{ht��E���D���E"O���CJ?f6��Q�̀�l�dy�"Ȏ�u!şc��$�WL��&�,�@"O�a5挠{���k�8	b�2�"O`��!��R��
 +�<���"OR�#�c�6ur����	<FP�X�"O��yqN�b ĝX"ɍ�>:,3�"O��[�ĿqYd	�V,�|3�"O����"W�S`��q�(�e$����"O��Ĕ�i�,Ke
��+���e"O�(QwB�~8���V㑪O���"O�S2,U%Hsh�`��&+i+$"O�q�"����H��DԂU����"Ox	h��Vos�(q⑈(�\p�"O�����E\H��D��E���*�"O"ach�+Ђ��ƎV�Gm�m��"OxȲ����r��c���V���9�"O��!��S.`�<�񉞜�d-��"O��cR��J����W��	l����`"O�!3��Z��IIB#ݑsn�٫B"O:��!@�CEl�0��_���"O~��4.ˣgr�0�S��`R��iu"O^��r,��(��ݠ�
�<wQ.p�"O&�:��آG�ȵ�Vc�'8n��"O����bP��Z�R�BK;` �|""O��z� ��]e�U�Ē�d�Ѝ�2"OR��?
�6���S�pNeI�"O���eI� �Ĉ�Ʀ[?4 ��"O�L�e�ۙ9lx���V<FX��"O � �/��V7$̉��3h�� S"OTA���S*�RTMѧ7�D�[1"On1(����PΪP2�����}��"O,$y!������]۪�C�"O$ ���8Q��J� �W*���"O<Y"!�M�f< ��D��7(�)�"O�����z��肁�ȣt�P��a"OX s��5l�X���������'dٱ�Ċ7��5���*:[l�
�'Kb�[[x����1�����'|�q�ժ��P��4z��@�� ��'�.8�ܳ-�P0��/>�bŃ�'�rA�5�о�ș���4:`�LZ�'���!,U�^��vN�����	�'�:{�n�e��5�vӵt����'�b,��i�,�Z|"��	���ԉ�'�[Fg�4c��J$�[�(��}�
�'jɲ%�C�7�A�&H��D�t:	�'6i�w	ô=�����Ił���'D
8�a�z2h���)S�5r���'Z>)�E'eD�9�Z42|�
�'���a��NdL)tF?!8`9��'qN@�E��r}�-TRt�+
�'�*�X�%��M�Ԭ#b�� 
�'���J6k³�fyw��:$±r
�'�(h��,������5"�(�'�n�Sbd�*b��:�G�=)�x�'�u8sa3a U�І���>���'A�5�E�(�<:�Dׂ�MP�'��4
�PcAsq"�o�6 ��'�P�b�@�|�TQ��Q�N`�'��k�Æ�Vo P�t���P@� ��� Ȱ��P|�Hqh�6K��5q "O�=!�!$
b �&�o�Z��"O����#	57t�y�B啄<Z!˒"O e;C/�Q5�)҆�+tu�v"O��Y��C�l�Z%&�~������៤�솰4�F����
���ks�'"�8L���ɒ�� �4s���Iǟ8ɠD��"|�۴Y�,��GG�$����� D�L�Ez2�v6mْ��]��xq3E=���S����U�p����
B�'S���?�L~�ߴ+�e�@�T4������9|>y���'��O?��	0��8w�Z�1�,�JUI�PI�	��HO��E��@��ɦ�S	�ak�as�唐mO2ܨ砦�(3���;(A�|��py�O1����x� (m讝k����h�s�AV�
��{��"fY(���1Of�4�f�K���U�8B�&�.=1pi2<���_�Q.౺���s�}�$ˑ�������F����6O��̊h�&)����?)�����O>7�@a�.��n�'��0k���Z����O��DʆBR�����.����Ƈ�"��'���I3�Z���y��ZilZ52�B���e,~]�3mИT��$i)O.9�s鑶?bX��v�i�!����B�F]8�P�͌ ��	��Pb~�8#�T�����@�g�R8�q���=�
3�O�>���[V>`�fmX�Lj7'�O����H>9UMʔǰ>�w�ڟ��Iz�Iڟ��I~}�E9qs��"�m�w4���=�~��'|�d�3?.n��G�>��%���!T����$��	�🤕''������k݊�s��8`�[�&ڻE�^�����ޫ�M#�y����A��UY�����т��$J�5K�/E	e2h"��'��X�"�"i�L�����ēu��>Y��@s�	dx,E)��'��h��M#���L����/H�D�Q1M�"7��O���?Y�b]?u�P��>H���t�_/Mm^Ih�G$��E��>i6	��?����B�>��Fc��4c� W.�M;*O���F�	G�&�i���Tq'M� >�� ;����f��r�T�w.��I�Xt���Sٖ����֙=ց��杼<Y��8��K�#=YB	��,��PZZ⪓�F��ӧ`}d����!bܘ�G�4|�#=�#�����	��M3���	YYl\�C�H1���Hg��yG0���@�S����dr����M��}��q�`� 1割�HO�Ө$�T@�4�MKխ�P��L��#c+d@�A?�q� �R��S���4��D���d�zF3f�Į���uh�><�v���	�WK�T�1�~���i>�8&��n�}�MX�N��y�
X�a�ؙL�\8o"2�4�S�iW�@�� OҒ^������f�z�[s��`@倯{��#&�i���X��?1W�i�2�s���/І����A�Z�དྷ��Ov�$<�O��f�	����tM���"������T^�<�D(��h�u��H;z���h˲r�>`�t�ٛ,�<AO>Yۓ!���  @�?   �  �    �  �&   �pA���d�Zv)C�'ll\�0BLz+� {�ɔo�J�H	��P~��#/�+$�^9��
���}0d�1��8c#���">c�M�V�8!��J���#z*�K��ӬI@��dS���ē�GR��"A�YAZ&$���'d|��'p����f���r����B?��za%Pa �{bC(�$� ��H鑀+ʨkaC��:�qO|H�q��O���8�D��j�A� ]��z��ʮDŘ��g�D<|b�X�bK!�i-u���=��@w!�B�!�d�'X]*��1�D�10ǊT�vt�
��O�)��%�x�a�H�=͜]��'�fl�0��%_���Q�.E~P����-�S��/R�"�S�ap!h��ϲw�ўdb6d��'��eΧ.��ѓsi�]:�q�@
u��<h�y�A}��|�}&��0dOӀBщ�o
�-%*�C�`4D�,�@��%F�HC3��J2،��1�J���O��H�����`�#�2�)��'��I @�A�C�^��e�/%��r�)ʉ�-�;&��T��N;$�ɑiC��?iҌ��v1O�k�2iM<�	@�MP���B�!BQACD� �\��d27,l���֍a�r�S�`�y�!�ՠdQH�1VbS	+�btX`H���4��	�36��0RAmZJeC��	�lo^C�	)"��q�Ĭ	����h��u�^��Ob}r�8ғ��'���E�.�&��qBW:x��	����:k�X ��2�I
[�&+�y��/<��H�ط�xhb��}�`�0_�e�`��dU�_��4�ю�V��r�?"Iт�NA+?�6���[H�1�EN�K.������ VD��'>��'("U���	U�*�v�д���t�� 䚴 �2	��/��o��L A�T��Y���~���=�؁�?��{�@ [�B���46�B����ױ6z~1���A^�^��8rd�E�]��$?E�&�Ze���A/L�5�9#U�5D����f	�f�h9�0~]��M4LO㟀��kٙ~��q�R�K(G�l'�1D�,�C����f��hG3m�t�g�)�	��HO�S.��$#Q 	#��m TJ7d�q�=����1�`q���͟�|zP�V \Ti�K�-&��A�L�3��I�mE�������O���'%���C�t\��b��1CUz��L<�#O�����O�(��#�]ڎ8 !�� �ē"�������&?�$>%���ʲw�R�����Z��K'c4�����	�5E6��׊ѥ/%������� �E{�O ��<1�*��q	�� ��?L��}�
�y2�'Z�ɿ��	!�IiP��G�K�'La�l�V94��'9xk�'��#�#hX	��	�4��hk�JRY��$�>��ěwX�l�P�-	�ș'�ԷT{<�{ǩˆ��'|4�[�S�g�	�<�f�H2j�6��$,�8Z��B�ɇ)�I:�M��~��,�s�7-��'"=ͧ�ē�J���+O�,,���C�"}v$���å������IV�&�~킆�Z�K:6�ɳ�E�7yZ49�B�5^.�9�wc���2A1F�txq��Da��s&��3ҕ��1B���%G�Zb��	b�u� D̟@��~�I͟��{�U*�ai钣*4^��#Hδ	�p�ȓk0I�'�A�n�6��	�":��=�i�R�l
��C��M󨟄p�)�`��m
pIM�{�*�Д�2��$}�]V�'6��pOJ�8�\��nQZ��p	�gN���g땺��	��&c��$��B$n�-i��d�'M����?��Oޭ B��Ze3�S�]��;6�O����OJ��?i�̾:jn�Wg[[v�G�?��hO���0Ǝm:��#)6 ��8f��A��O��� ��<��$��B&Kx�M��#³Z-:����W��qO���ŋ�N�g��+�v��4�C.b�H���K6�BB䉦c��<H`%ӇW:(-��̓�+�tb�E{��df�9}/��4��h����
	�'�(���,��-�7dL�Fp�Q��)���1��`�x���T ń�~rh[�ܸ'�>7� ���Ҵ'v\�J֎	�kb\̸� k8��d�9d�fXka�ܛ	L�rQd�F�!򄌍?�Z! �a�a����χ,��Ѕ�	$�<�GeF�(9���E9:�B䉈k@Y���	<�����E���	Vyb�'�ꍱ`L��0�����'T�Ze��O�6��t�qO؄quKQ:��y��8�wǝ:�![�M�gm�̆ȓNE����ㆺ]�
�Bv��9d�Ȇȓ������L��Y�J�'����'V�hi�����)bdJe�Т㓯�
Fv�(�a��L^�$!d��.4Gx��ɽ}2���A������E�51T�� Z�6��O�x�{R'm�SFQ*=*d#E�][^��2L�3 �B�	�p�*8���B�{��p�W�&K����.�	Y�F����4%��Hd�ԇ��B�I;;ݢ90C�D8͸��t�
��"<����?�QPo]�ge�x"P�G!�Ĭ�qE�_�'�P�{�G��?��҉�W�^8�s�Ĵ,����fܓ���E��xR���7�>�+��@~����uJG��y�a�4_Ģ�����9!gj�ԡJ��'Hўb>���Z�B���LŔ&@1sL*D� �E/T�emT0�Q�P�g������[���i4�	`�Z�X��T28�;g�n��	%iY��j��S�������n�t��%�J3������6[��⬗���,�ǱPX�e_Xr$�',� #aٮS�yq�
�XJP=��$/<O�L�ț5h���A!U�)7
�۱"O��㣃Lf1�
�/H�76O�˓�hO �Ot͒t���"��1�0�-8�0���V��mڼsL��<��+������pV3M��$��H�!�$��w��qz�h������K�!�DX K���E 7r_<|ZV�P�.��C�[*����`��5k|�+a��(����;�$ȵ1���:r�Ы+h�("m����~�J��?��NV�=R8��g%J2}��4�	l�|*p㞬I��4f�q�0��F��/j��Q��5�y�	/��X��\;6�Đ�3$�$�0=���`��F���b
$!�陃�5�y2�Հ&��\8e'Ѳ|���`��Ox�=�O������ک�\����i���R���#G�qO ���e������!�H�Є2Fqn�=9�#'����':�Xc"�8U4���4�7K�����'����d ݒM��dO	V�u��y"�)��pښ�b@�,~��` V��LB䉃���%�rޚ�jw�-E{ʟn⟄b�F(�����-T�]BA��+q���&�Gܓ�MG�B9��Q(��R!2_8IIW�#LV�D�c-]W��s��äA� tJ7�ѤB��3��0D�Q����q�`ؔ B�X��l��/���<�ǅ	�<0`�L�y;:�,��ȓR�Щ�����~�.��G�Զ^�����$6|O�)E������,�R�v���T��mZ'c0<�<y�:���'��(Ƅu#�x����/ !��lG�}2�(V!∳7�ܴv	!�D]�;��u�� ](&�Vi
 `FC�ɎA���"bF��e�G�̈6vd��"��n����	�"O�����D9%�~��V��?q�I9FO6����u�����M�_E����Q��doۗ�h�pa���"a��A�⚴�yd{�%��Bж2�Q��(�0=	�m܆>��bڹ
� �A����y��5��Y�''ɠb:
_5�OУ=�O*:@H1'�i��%ku� Up���g%ғ+�Yc��	�Z fD�V�Ig�X��"O� &��!'G�_I��H��ޅe6����"O"��bΏ�:�� �4r�g"O�Q 2�Ll:��E��l2d���"O6����i������$��,��"O4Ȉ��ݮ2�P�R��/�.q��O�h�q�)�'j(���*ɴk8,�B��:v����O$q��K:Δ(9�	��AȶU�����WKM�"�̹`� t@"�ȓ|���� �� #d���{����K�f��aJ!O����B�t�t��ȓv����H*�`2��:�r��O�:��'w@�Ѷɇ-�&i�����=4.��'��"SM�<�t kC� 0FR ��'\����bS�'#����LF1m�A
�'��u�e�ÀG0m��ȖWG����'�&�f/@YJ�3$��&SJl�	�md���	�+�ɣ����8��oѯ�C䉦J�a��U5QFƈ� O=|�B�I�mn�S��-;��
1_jB�	v�8�Qę�`��H�̓�9�C�ɪ����ּ���@�0�rC�	�$1�ŊNeVd{ց����>!�-�n�O8��R�9ya��+"J֐	��I�'�TP�.�R��y� �*|"ԫ�'�dQʰ�K�|��X����*b&8�*�'*��Ó7Ui4h����aϒL��'̎Q��J݄C��������`�	�'�6S&��D����B���#�'��Mۍ��MTX�B&�Q�o��,�u��\�nB䉱k'~�c��̬
U�G	�B�I�O�N1�D�c4��!��&��#<)ϓZ.ڕ��C�*P<�Y�ʝ �I��K �L�$�ru6-1b��:gb��I���In�'K��O耳�ҩL�����؟N��ܰ�O�`*��;?1O�`�ݴw�|�On�)��_=,��Qa��1�j���"O���$"�~,´b�-)���"O.� �c�.l��`a7EW�/n�H!-4�y�1�b=��̌-Q!4�	��5|O�&���7+��@�J�P��/�rr��9�Ix�'
ţ&��O�i36"U���ʱ�L$i���>)rlH�H-p��<A�ÉY�?Q�F5#�"йa��\�Á�6*�B��5eg���-��4T��7�N)�&���-�	q��Q
G �|�D�"EO!y��C䉐-�<̛U���BTӦ�˗H��P���?�H�iK�p����E�D�.�0�Ll�'�R�!��#�2L��IҜ@ l�&��{gv%ڐ��8��b�"7.G�q��'��I�m�3��aYr�^�Tۘ���'�2�:�����x�.H�S��� �y��)��q�j���D�/�ZxaQ8"��B�Gk��@�Ƈ�� P`��"[�Gz�X>5ۉB�yJa��� ��^1��LQ��?��GˉF71Oڤ���N:���a�&�()&�y��E�`�1s@�ޜi�rn_)	6䑊�I�5~�(]����yo�������M��t��]�0C�<�O�����5JI\��#L�	x=^� �<�!��ԼO��H�gK�mY�\�t�X�C�⇮>���IV̓)�q:�ʓ������ⓙvi���Ma�8�
KK̓Fa�7M
^�'--�|@�)M3Q��y�%��d�� �ȓt`B���n�h.�t��g�z܇����4a��J@"c��#[;����'h`P��It $�����$S���ߓz$�'w<@�W�MV&�,B_D���B�I�n��!�	����gH�89E���)O�'u� lZ45�1O 駞��O[�O�F�KQa��0�-��y
� 
yJ2,\�e�t��t�� N�$࠱�'��O&�!��ʓ$ �z�Pc�l�Q�"O������b��Ա�ڿ�F䱔�D�H���i֮iW@�� `��^�4L���=��/S1O* ��O��p
����p`<��c��,��D���$ׅQ0ȸ���L>Ar��>mˌ�	Տ��II�"n�{�<�7蛡?�֜�1�B*�*�E�z̓�hO1��AA�eX�~�(�f_5Sq���"O�M��t�h���_2|a���V)<ғ���r�f����B�"t,I��H[�9 ���l��mӍy�Fg�Oj�����<.��ز1��rQl��g�؈T���L<P�D���%��j����/Zb��3��+3��>*c��a��� :��Ex��'F���Тɂ|A�P@&ťt��I��'��d"���*���� mk�����X��ɀ�HO�c��pQML|�V5y��~�Hr�)��ܰ6�	�w�c���v�i�zp'���t�X�m����)@�Y��0IG#(D���b�N0�H���;F${"�'D�e��O���P�`C��0"7ŏnh<����� �A��jd�EʀZ��@�H>q@��NJ�r`�-�|�B�L���hO��ڑ�Yԟt;���
 ��9اc7_��ya5�"}rL�Ӧ�9�X1$#�O�QkDHS�#b�픮�4��'TXKAA�	\�u��h�z�)�ӓ��'8��l�}iJ5�G)Tr����'Q8�����B��C�'�W� Z��5�S��߫��5+Ѣ̠3�\��*�x�"=	# �1+1O�9��w�=ZX!n!�t��5=�N�B���'����S�g�	�#�� y�eB�V��Kڍ�C�.x �@�͜5!�R:e=z�b�F{���,H8A�h������c�+�.�yr%5f�� !�	 b�p�4]V���O� �,���3h�@�����9����c��O��x�p�Z��|�-�z�M��m��M��dl�}�w�K�����(.���i	[�@��1D�X[��JnJ1�䄀y��A*��<y�TLATLy�ƒ����`��M�<�dO֪@�ڀ(`Nߙ'7<����Ɵt�Ol9Ezr6�͒h�F�J�O����7�H( �d 
���S�ɪt�'m��կ!���`�A:'�t���'Ѥ�QoNi/����%�2%1�L�
�'F�0x��wp^l�R=H�P�O�mS	�m	�*�t��蘒�'�ܒO�ey��H2>���u)_�Y:�s��]�'�E�v��OF͠B��#}� ��Eu�	��>� �.u���<y���Q�S���P3,/JV��
䬍7*}�B�I1z;~�5���b���Ya�� ����$7�I���u��&?��) �O�~r�C�ɂv䚱1�f�y�,9�1L�-vZ�`����?�p�Gďq��X�P���G��0 ��Q�'���#�ɡ��i�r��$�2��.It��&/2xc�0�V��`3q��'T|���ٱ,�̸QB�,0R愐	�'����V��%� j	�)�y��)�S<2�KJ�K�@�k �1!���S�"O��u)�)C\ OA�)���b7ғ��JT��r�ɩ‏�M@�5�ć�%qέ�ɧ*�e#�y�Ϟ�����V
ܝ�`�Οy�`���Q5x�nY{1�'��2��7m�,��ʙ7� ` �'��	cDZ�c���ڷ��6�^Q����4<OX�
Յ��K�<k2�X���B�"O�a��&��<����q�����'s��ߑ���<��	z�"��4q�,�e?� ��/Zt�<�Ab�\D�H>�sG@���AS�"Js�P�re(�a�<a�-X� ���p�݅M�м�S�\�<� ��ї+���p�@ηAu -rs�74��E�gP� ����H?�i[0�+|OV�&��)Tcڛ�d��@h.d���*����HOԝc&���#CǊ�2-ι{d�P!K��`a*�	�.1O�\�B���#�njb�)q�E� � �q�ұ�y�=jAp�[7e[? ���qfcҟ�0=����-a�BUqpg����IO��yR�R�H"����]7
)����I<��'�#=�O���`l!!�PXˤ�٤y��d1��	9��堎y�!��|r'�q�\�#ǐ<��ݣҺ��c�Z�mU�^�q��'�����m0��g�V��1�'�r��AT�@JUk��� R�F�y��)�>S]��T(D�{.b8r�ѻzzHC�k�ũ�@�3>D"!����
��Fz�X>%y�2�R�LMcE�@�� #��	�.���%��8|{� y�	�g�t�s�_$�|$xׇ��=f��r�L�{6� I���?Y!��i���d �L<�`%�� q @�M�mfP���E݂9>�J���4�ߕU0
��~&��iR�<G8�<�E�ڥ[(B�0��?��O^��e����ɣX�S�.D?!�Xh�0�ܩ��C��n:�pdjݹ;N,3�[�7����<�F��r��Rv�'w�I�Y�YA�gҖ��m�4�0T�jİd��:~>�Fx
�Ҧ�IF�>�1hߝ�u('!	�%�A+N$b�!{��_��R�fW9)�,���_{�<[�h�#h�\�:F�RS�L�R&�@�E�Z���3Wj���d�("�B�ۗ��m�l�bD�>n0��ٵ�'��d�-�>�����=?�e����>V7���ɤ��!���q�/۩=[~bu�^�"~���=A��[��?��{b�H��x��[ V'�	3��U�~�$�~U���7m����'�T-�M~�$��]���׮�<b�d�J5�i�<�d!Q:X�Dk!�5���$#�c��H�?��c�;�@X�&�2�(=��"SZ�<�R�@G �qBͶ~7`��W��W���P#�=���nJ�+D��'R����I�n�(��yR�|"C��?���ŭY0	�3`�Z���'��8`�Zv�g�(� ��4�nE��e·T��C�
8�5����5�P�+U09jb�TD{���F5%*9��ϚkM�*eǞ��yR�Ω5��(133@�賤#(�����O��㟈�7D�d�J�ʀf˽T�X�HU��O�1��A�T̓a��1F���ױ,%���×�D�Z� e�K��\�P�B,��?��v���1a�$E�;q^\B�	?3p�������W����fG�..��"<qϓ{����Po��6�)�ƃ�-�`��ȓ:�0�D��Eei�f2g�)�ɞ��$�G�'���O>A����S�l8��U�TL�@9��O���f+�cS1O��J޴ ��Of�JB�9n$��ZD+!z$�89�"O���!� ���j� X	�a"O$���|d�m�UIM81�\�3��-4�H���
R�΁s��u�D�+|O�%��#�:�:3d�1 ��,4��b�'�
��%�O�5���`(ö$�53}����>醍˥k��T�<	�Z�_�2MYr�LI�t��ԂC9bC䉐SK����L�utpe�ίZ{J���'�IB��r���)ςR���%}hB䉴6Iؙ!d,�r 0!�EL���@b���?�c�KP�!�ީI��G�4$2�[�ANJ�' ��c�7�ɌF �i�� Z�!Y��h�܀��Ó���c����q��'���e"�v�yH�,�=k��E`�'���hP��xJeȮ5�s��� ^1O��=�|���,,20S��e�<A贄�K�<a6��D�Ƽе�ǯ/�9���Ɇ�HO.�'E�Oj��p��SՄ3}�:�0OR���ϿR] 4  �    b  z  >  �  �$  +  c,   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�H�!xn���G*W�(:h�.|&�t�BfE�C�V����5��8b��M�5P>D���@$K���x���1Hm�� ֡mD8�3�̕�Il2�"�JMz�8-�t99��'d5���!"ӫylhQsϒ�UT��VJ7Q&��&݅tΨA#�7z]Ҝ˴�USX�\8��!s��L�;u^"�z��9D�D�ҡ��[�z�{U���Й���*D�|!�*eZ�h7��K򺭁�*D�H�� z�.�ك/%��qu�:D���߅Mu� zBb�,5�f����5D��ڵ���?�i�d�R?R~�覬8D���RF�  hyI&h��D����&8D�P�gmܩS�d��wቀ`v!0w&8D�ܐu�lR���W+6�p��Sj2D������~(I���;�`5�#1D�h�ŇOB�t����Q�y>!05f=D��+!b;��)��p�X�(6�;D�8kC�|���^�gHP��6�<D��ʳn��v�Ȕ�-�IP=� <D��
�����P$�9v��!���y�B�9�~���,�zi�I �nފ�y����w^iZ�n[w 9f@H��y��Z3;+$L�RmT�7���h� 8�y¨�IFܳ��V8��&�ɹ�y"d�>xRLɋ�ˑ�Wj�ƌ���yi�$�����N��\�b������yr$�twj��0*e��Ā*	�'lp����=A��������=����'[ZԒ����􅛱��&;h��'-�@��Ш�D��)F�H9����'�@}���0c8L�F�
�A���	�'u��@K:ɀ��AF K�x��'by �,S��>$q�FX:�&x+�'�:�"��Rx�S��R.,�~���'�l��e�S�=���+��ܒ�'~v��锆P`�+��[ze��ɲ����w�^!A�!��lU�<��5��@x%�DY�T�ă>xa{RD"8 �����6+Tm���ӈO
hC��7!�b����p;a��u,��HaZ� �3�"\I�õ�ybBL:ւ�;i�<>*�Caÿ�yb)��s����᧚T��:bFD�MG��� c@� ���.����B"�
�y�$�^qp��N98�L({p(�=R��Y���M+�EO�E�E�?5��}�	4I�,X�k�U���5���0?A�, I�%�+x�|d-YC�����,Z���I�7p�Г7�'00Kg��>|+@�g�իE\کC���F���Ӆk4���{��C+U�^w��!œ[Qb� gb
2R4�2
�'�XXU�Úr�2D)���_N|��'E��(�-K�B^q���Ϫ��X �t�OH����Ip\�p	�m�)
�'�^���m��1���FL��D:�M�G�)+�F8ٴv�)9�L�i���7��'�d�j�"<���p5�ذdjΑ����I;'�]-���D@��Kl�C�!Bk�e`�旫nD�����F*D[a{R���ԥ����RN �k�ռ��O�}������PU��Qmb��U��uJ7HUC!MĴ[�!��L���y"Ƀ�#f:�I��=���R��o?1�ED�/lA�7耆j�����E���#}���ə��PA��|�n���U�<�A_8D!{�n�_�P��A.�&NPt��QE���PxHE�Ο��>��	�<g�0K��~���Ug���s��m�fʱ�(+�eiU␬8�r�`а<�Ή��fS�ve�ɻ�t ��I��V�0�$ҙC�D�F|���.��8�SӚ;�D;ql�8�M����P�e�����@/C4��Ņ��0e�$�E�r��D�[�7^���j�ܔ(�Jðm�>�y�@	+�eo:�'M �aQ6�J�[���c���.D2}��l��UЇ�͠_�f[2���z��	��LP]�ZoڼB�x�WK&���i�{d��#�%��Zs���|Q�0��I�:�"�5� ,��*Y	�z�Q���?x&Dz��� ~���2��	E����I�R��i����!
,ƉQ��/�4#>iSnW&mS|:F��(*�4��!������fhǯ"E��U��dM#�"C�ɟ'9^)��'�!�ؙ��X^牒x=��p��)a��Q��؏y�7�Ӽ:�@Cn[�����&�(��B�Ɂ�Fd��B�{w��z��˅���oL�o7�F��Pq�'R�d�6���5v�ѣ��ϿaT*�j�����@����|�D���P���<�T���Z� Q�B����xr�ēh\ yc�_؞p�'!�2�+�/P?`
���7����`Q��A�x�HI�C�|�oz�ey�2:%B(��(���(�l D�zP`F~���� <��H��n+D�� P8l�$�0�΂�s��`3Ŏ7D�XEӮ3X�	��d%��L��*6D�
�^�S�b�r�E��`�)�t�5D���jW1%�0	W$L�>��Emo/D�PQ�
5F}�; �����`/D�Xx�<���BfP���#+D��z��D�4>�B3�G�,��6D� �*�,08R9y5D 1{&H�@!D�����8T�z��lܥM$�y��.D��#��R#�̛����w��c�'D�T��:XQ���5}�*���:D��I�LǓB0j<�sU*���R��9D�x���U�<\Pvϖ�0b��J�M3D�(r拖=FLAI�*7*�x	I�2D�@�5��2Q0)�;ydc��>D�A�t�܀ƌ��o�ɉ�:D�Ԉd@�i�.83
[�Ӟ08��2D�$KO�(()�eڵ*�i.~�!�$х<��)��.�<9�d�f(�,u�!�$O�6��2%"��r�:8���;B1!�d�&j�2N##��\�-��!�ޅ9������;��V�D�F!�DQ0���C�q�j�4lϤ]a{"&I����'Hػ#��{@�bl�4��/���(�g��l���[�fI�<���K�&�H0���жA���ʔ�
�  ���
�!��1s�-����cԕ�*�4�>p7�"��B�@���~&�� f�ܗ:���#B�H�(�PK,4��7�^�~�eK�!�/hZ��*�lG�1��	�H�����$̹j+pX����6HN���Ҝy��y���v�N���¼9>���E����Ɗ�[�pbS��!��חoDZuF�ɚ?��*ᦀ�$q1O�(宐�d�~|�B�%ڧw!l�(�aArg,�����'L���ȓ10����?d��E�E0^MW��_8���It?��b*��D-Lr$�  *�08V<��⟴M��Lr��Y W-H#��#�ʶ'�T��Dk��5�rԀ0��8~R�l��	�S�C��*2� �1�V�z�F����d1Pk
�hu��`�o�tB�%(	���#*߿g�,���R�d, F@��%uN����sYJe&�����63�Jd !E� ���|�Q튆Ӕ�q�N7	�(��5��z�<����[�X1��L�*�q6ǌ�`��a�hL�	�!����O�Ei��K5_'�\�� ?7l���'8l��D�3/����C��,�E�ԥR�g��8�ff�.|���0$&@4��z�㟪K|�I�ADD�+��W&ޮ��OT\�7F
/b�"4Z�h]�rqv���Gť2�rxY3I��x(`��'-�>��,�ȓ@��)P��ec���S&>��'�@Tѓ���N��T&��&DD��ר.����`�9O|���B��y���SU<-�0E������C�nn� :Q�ÂH�T��'���!�|�=�iB�F/�!�@������.	����+&����"d�T$)#�ܛr�5�&�B�?�\ @�EU�r̼kߓR&^�kA#Y?0�@��<�=��I+ZI:9��!O$:���Aɟ���(�.5I��[	�9��*=D��Id4�X)��$|F�e�5�x�Y��KE�w	l�~� �Hy�D�7w��,ッ=@�HM�"ONas����P�e��.�C3�g1ȉ�,OR��S��]b�np�	�gi�#��͙SI�I��1� �1D�@��_�Nx�r�աA��C��<9�>�� @������<\�8%�Ī@�c2��'N
2YEa{r�P&x�x.�8�ӕ*KN��R05���R�#<\������=�d!��<_��0�
��Re�$�E}��@�T�N,%)2u����ğ����6"(@��<D�O(D�x Ab�}�@����ۊ`������9��˪ L������'R�V0��S�W��!h�O� *�� �g%�@��B�I�\m�$�O�=/���y��ƻ(`~���NX>qd���O�D��3?�Db�9@�\�J�c�-;�����g^D�<��G��P�	cmE��|���A\ݦ)R⟶`ᬬ
0h�/�0=��/ T&���e�1|~���§Nc؞�8��>p���k�O@�8Ȫ�Q�u�[��4(����'���P�/����[��^'����}�Y�ka���RK�\�,���ZM�0I`@�NVTd���{�<�p��GlZ#�č�=�� PL��1y���u2J�j�'�#}�'�l hv��^�ހ�Ёզd3"��'ɬH+7��n�B����fc����2J93��4i�ij2�'�R�x�	\l��y��J�
QE	Ó`�aq���4�V��� Z�2�z=KGϐ�=jpp�N/B��ڧ`����x"ʐC��s��I��)��
T����Kd�Q$i�"�D�FkX�7���?�Z��ȡ (H)㨑�T"�:U�#D�P�`U�kR�<*����FA�i�!�V4�"m݃��{�g4_�>�O�܃�K�4T��:RA5A %:&
O�@�m
�QH�%G_*t�J���:P���L���� D���0=qEH·K�>��Ņ?w��ЊФ�}X�|�#�+?n6���Y?;.����Y6h��MB�vx���T$߄�y���CR@
�|�����%��ēYx�DkWA[h�ఱvjX*�(�~(*c��[��5� r���q�"O6h�� ��+�S�5Z �auk�/��8:�j�<$��M����@/K��1��-�Ƚ���>.!�[S�j�+fK��q��-@�FT�@��3�V�"6���+|O.�8�HY�I��ձu`Њ91�<�r�'6X5/V�'���&d�C(�\0#4��J�!�R,qL�R����@�6�ʩc/�P;q�E�Ob����d�#+�ޤc��Ά+�:���'�`BDI1o�xahM�0E��'),Z�Lԩ^�@)A��ߒ�U	�'��4�2%��>4���7\Az���'o���F�K�"M�A��M����'���[��ߞpnx) '�I��`�'�� �Q@ʅcզ�T��:o�\��'��y��+�T+�j_6`"�{�'�NI��i�DA�2	C�;���'�d)CVN݁t��pc"F���D��'R��sˁ��ㅨO#	�]y�'3 ��7+i��esGI9v�`�'�젨%̃~䡲3�	{��C�'n$I�W��:~& ���T�=�� ��'�T�zs.-5�<��3�R�K�'^�<j�H��B�$�r#ч%� (I�'@N\���[�z��T`�ə)�)��'�-�EN�.%��5'	�	W�1��'c&�t
ɡF�!�&5�	�'��U��O�J��X6k�&X��'W��sH��n���$J�$ ���+��YU��VN%�L�hЊ��ȓy���;�њo��<�� ���]��y�i�3��2hµ9���\fn@��5��X Q��RH���˔�~�F!�� �x ==� 4��hF���ȓL T����*��9���*� P��S�? @���E�GN�h�jеa$��3"O$H�"��.U2u�!�\�K�NiZ3"OX���ԓ:ZzY�7���L���"Ox�jB K2_ւ�8��̇g��X�"O��h�e�Pj��;�aH�V���"O0�[E�W���К��ϙ0<p)w"O����3�< ԡ�V�����"O�I���R!IZ��[0'V�Ep�L��"O"������A�bh��B�"U�UG(ʺ�Z��*�vX��0R	щ}���S�-WӦ��j#D���d!Y6-��,�����|Mi��"D�Ը5+ Wbd�`͞�`I:��+D�t��b�56��R��]�X�B]��)D��㤢�'#�#�A��s
Ջ��'D�8�bQ��v C�ѵv��i��&D��Z%d�??�R0y�.͎I59�P�.D��'ϛ�R��	��M�4��F� D�dI�m#~�譨*�\>ؚ&�=D��a��[!OQrT���tc&��:D�H���D�j`���2Q![��[��6D�lsL��@ɚ��T�k���i2D�h���%.mN9�H� P�m�բ#D� Q��%=�ʡ�ք� j��$�L/D�H�pJ�.|c҈j2�L$%x���)-D��[��D4��@'�I �X�ȗ-D����&Pla���S�T�R�Ia*D��35��3f������+<�v��W�*D�$+��Ƚe,Xc���a�&���=D�|r��TU@pB3'���怲s�6D��16��')(^,:"��`����3D��7j��>	(�F"� ��83�1D��k�U�X���QW��)"V�� k"D�Hz��#r���!�B<P��� !D�� e��	4�:�1��^=j�(<D����	�(��ܒ�L��rC���F�;D�dX���Z߶�Ӆ��i��hJ#�+D�Ԙs�O� 5A1U_�!�"�(D�`Q!M¨��1�Pŏ�A5F̡��:D�h9���P�������/�X4i�+D��2���'���hJD��D�<#,�����3K�T�5��I[f�<)�ʛ?�pP��Q�����EP}�<4Ajpx]{�,C����K�f�z�<��M��~�b@f�"�h�3DM�u�<q1���S�j���fU-��$#�t�<����:%{�AęaEH8C�]F�<����IB!*ZS���LB�<�e�`4R]h#��:�!J��E�<1��:%H�1��?-AYP��@�<�W*_,>�z��%��y�J_E�<��-��G1μ��|�A-�J�<�*�'�"���o� hY��9)KD�<�$���N���%������`A�j�<I �R���qp���D0`%�D�f�<�c��>K~X���D>ϠP�ef�d�<y�M ������H$� s��j�<��)�htx ��l=:{��
��k�<�d%�1.dT"�._>�կ�B�<ɵ	�wV@�I&D(QM.��G{�<ylM%ھ���	<(��H���Q�<��f�h���bؼ����N�<�F!Q���`�HQ�4|�E�P	S�<Q�5�-��a	�8#V�%�VM�<�tN�i9�ĸ�ႁ,�"5��B�K�<� �@�� �k|T��O�D��"ON<�ƌ�6�����.�oƌX�"O�evHɳ5�pA��$L�X��`"O�`�?E��Pk'�h�^9��"O����"�;ȩ�V�P�.:�U�V"O��QD��2��U�!oQ�)0D�%"O���ݹ����+3���"O��� L��Ze��Q+&̉v"O΍����s��q�r/�S22��"O�T���2g�4i��MHH�"O|ؒ4��s������>]J�"O��g�U��26'�1u�
4��"O�|1��#x�b�s�/D/v�!	�"Oz�JA�S��y�� ?G:t��q"O(���+K�mՔ�3ፚNzvi�a"O�-PE���4XW�Y0$`��P"O� ���VTZ��2w2�)7"Od!I`j͈
k�0^mj,
�"O�y���D����Ca��	l�*Q�"O�e�㌍�6,��H���9��kA"O4�Q� p!�h[Ķ��J�"O��U	�#��aK�ԿI�T�p�"OV`��H�M�&%#E�R�-WVp��"Oʘ1�L�^����ϐ�03&�3�"O�ᢧ/L�c����-C�W����"Oj�����pM�'��7QR��"Ol����ͳ$p�y�"��Op��0"OT���͘��~�[��!'�lHc"OpE9���x�P�3�+co���0"O�xz��L2�|�^<Q�:q"O�t���#4��!If��Q2]�p"O�� �*�l���ϲ\��[!"OlG��u��� qGY�u��"O1x��ͯI�����M֐q"O�w���{�l�q�āGPN�"OJiʆ�ę\>āӲE�#I�1@�"O��PD,S�\.�)v��`
��Jq"O*8aUE%/<,ͪv�	+T�h��"O�	��LщXo�x�H #fwxjq"Oly۰N	�F@�!cG�4 p�T��"O�|
�C@>	_HB��X Yj,��"On9D�Ȗhٶ���$u�Q��"O~ѳ� �)��yG]u����"O�mRG��69
^� �M
�a�b�à"O(����p#��RmF����Q2"Of���5��Z4��E����$"Or�{tgԯ^}�L�B���j��%ɡ"O�4���Wq��2+C��<�A"O��q��΢:�B��thCp�rH��"OzD�#��B�0<�!�R�px�e��"O�S$˰pT����5a�<c�"O�iCT,�/�R���K�R���Q"O:��#D���E�t���3�|�t"OT�e��Gr���CK�	��ݘ�"O ����=Z�CT��*�t�iE"OR��UGS�F��b��9>���Y"O@�{�h�</��$"�(��./p��*O����o��_ZLX�'؞>T��'�� ��!��8��E�/m��q�'�r�IbRZ u�F�/`h�`(	�'�X� �ϝ�C�F�`�������'/�����ސA��l�d�<J�
���'S�M1�g�a��
t�Um�#
�'S,A� �X��+#g$N���� X�!��7uaBh:DO7P�b�"O�A�0��A� ��eaV'{5�4��"O(���2d>X-b�F@W�T�qv"Od���ƀ&y`=K���IXt�p&"O�@b��5�rT�u�.��ѷ"OR�Y�c7^�F��Ċ�_����"O$$�1K�xk�H`4�Љ�Mp""O]�"H��=W�4ӵj[�_\t�w"O��V'>'ne�jD�S�)ѧ"O:YrC"���܄��Ɇ�gQ�	��"O���bm�+����(֊l�Ve[�"O¡h�/K,Qi���񡛩yي0�7"O~}eB�.Ql,Ġu�-���F"O���%eE9\?j�)0kU�K�h�+�"O�R���p��,p�C�qjJ�# "O�`����Ec�r%	��I�<q!�E-J���l��UТH�'C�G�<���B�/�h�S���9n�4)�V���<Y���3)Hb��g��qi𥲴!��<��͍+lŶ`�B��h;Ҥ��Bx�<�2W�'`�1�/O�mi��a�@\�<1��_
W#�����+\U�j��[^�<��/�p�f��R�Þ,P��f�^�<�F_Rm��3P�:��=rr%^�<�re�C����`�2UA�Q�<)��P�j#��q�Ɔ&6K�Z�nB�	��̅ �F�z�P4�&.޲IhB䉬 l4̚vD1X8���Q,$�B�	$�0�I���RZ
�9gB�1�B�I+��IY�,�s��})5��=Q+B�I�D���I2����J�_���C�I4@ܹ!R�<h�Q1b�ܡJ�C��'&Č���ޔ94Č��D�]�xC�	>v�D���W�&����3�)#$�C�	�l��x8aꙋ$�d!�S�:&�vC�ɧLn�i���jd�)���F�BC��R�L�� !F��<wC�Ɂxm,Dp���.�J9밈��Z�!�dK��,r���%tt�0�9t�!��ԜqA���ygDH�e�q!��F>0�j�'>@���.Jm!��\%�U�H��N%�m�`Oˇ`Z!�	���8�Zu�N=RT!�וshA�����7��0l��	�!�#T8`1f�-	-`�I
J�!򄚣c�r�r�CĜh���3c�	O�!��L.x;~�KS!��]XZi@��Y8Qd!�dʰ)���	�ݭX=)#�傠xU!�
*c��}����_V�t)$�1(8!�d��N�,���)i��� ��+!򄇳j:
�c��K!b��,B�@�E�!�G�#� ���ś�aBf���.��!�����=X�ƞ^4������U���J0��ME#M�>"��6�D?�y���x���3v��1(Q����Ʌ'�y��A�,�Z�3�V%$�\]�G��y"%�=�H��G�#��r �y2�G=y��@#�%�Rg�Ey1�Q+�y�fϮhH��˲kU �,���y���b=�,2��N?<H#��ޗ�y"�,>[^���A�=��q��X�y���h@��a��/�֝I7O�:�yB�� '�PCM��!��� D��y�ʵ�����?K01��b��y
� B%1����H䴱�t�]�@4���"O"Q�� )b�L��+�S���"O�I���:�����IS��L���"Ov�[�͎Z�Hܪ�ɜ9�^`)V"O��1"U-h  Qk�N�Ą��"O����^�v��d������"O�mBUh[�i��3@��&��L�R"O^�y��� G*¡z��3hh5k�"O��0�d� �D��E ��z���TJ�<�C�s*؊�$��1ж��Y�<���Y�k��m��!ջ�5:&j�t�<�&	Ĳ;)�	iDA^�\� ��c�m�<�Ҹ��R��˂{w�xb6mD�<��O� 
  ��   �  N  �  i   .  �;  _I  �V  �d  �q  �}  (�  �  ��  8�  {�  ΰ  �  [�  ��  ��  h�  ��  Z�  ��  /�  ��  ��  Y�  � �	 j  � �# - �5 �; �C �K DS �Y �_ �c  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C��'9�@2@��ՠ`�G��,i�_Z{!���[&�p�K@$&1���b�?4T!�]�S`d��aB&/ʘp%,�*@!�D�"h$���ԙa��K��!��S���ۅ}���bB��o�!���?v��]��Ǘa�N�+L�g�!�D;�:)����Q�Y:Q*:P !�$�yAP ��Q�K M8�I�t!�d��s�FѩdA�PrxLa)Z��!�Z(RvБR����wY�B��T�!�߬ACby8���T��tfH
M�!�W�`���)�==*��9�/D�aK!�d�o�ڵ,�1D�""n����'�X�{I�jG�%�&H?e�x9(�����(V8'l�A+���Z�!�=)��a�	�.^d�qE$��HH!�$�)R�Jy�Ӎ�&q���ץ.6���~|�ծ�YвP	��$֐��$��T�g�Џ!�� I�F�F�z)�ȓi���j!��.w�TX2����@��y��'�0�Fi��n]����- �#��ē)����ϱR�
!8�j�>A���ȓ.Ŷ�0�K$W��X�+]2`�@�ȓ^Z��I� r�Xƥ�2~BЅȓ.x*$�0f���ָ���o�<���
TtT�H%$yUnTSu�V�<I��-"���d�P�LAٺ�*�T�<�ad���Qpa�[�� �e_O�<�E�ѨU�R���F�a4�LH�<�#��:�`��ĕ�Z��� J�',a�ԠÅ99���TLF�Q���S�M� �y"����*�b��\P����(�y
� &�c�Y�W2���C+[�n> ���"O``��b���`�\��
y3"O*E��%�+�,DG� {^���"O�L��l�H�P����;YL�|�"OV��Fm�~wtq�1  ^���Ip^a����m��S��E�
pec���y�+�a<���A�H�vML�K�+�8�M����s�\�q��13�؁钫�_����5"O, �#L%D.F�*N=yD���"O�t9�/\�8BL�2�V�*P�'���0!K"-jE�_�Q�(�'�B9!�$[</Dq2V!Ҟ-��)��.)D!�ɖ5m �8��G^I�Xya��;s!�".�&Sf��#���@�ސ"!�$�.gg�UxU�/F�~�
LՁl�!�UX���(�(P�Ŗ;l��'�r��7���S� >{�V�#�˼F������Ob�ɶ}����� �(��GJ)S4C�I9���H�h����;��H�n*�B�ɟ{~^L���q�JR��?<�C�		?��U.H�RB�`b�C�T3�C�	hH����_�u`��to��r�xC�I+�!�K��\�<M��䒚"�`C�I"/�,D�F�3�H����}��B��
��`�pA��6�F#)@4�B䉀b`r�w�N�7^y��]�U�VB�I� ����	�<aF�R��ܽ=�0B䉘C�4#E�H4_�H�+����B��;��҄�v�~�B��pB�ɋ��2L@">v@�!O,e�\B�I�\���!ЅE�X^DpC�B�1'��3���q�,�C� E�,|�C��8�!��G!��!	`�N1Q@�C䉆t��1�J�#t_	���Q�V]C�I�/rTURd��/4R�!vJʍ5nC�	)l�
H����x�Td�G�<*��B�	$]� 9-ϫ���T �1��B�I��FC�i�,P:X�āF98�hC�;Ol�#���(�" zA��4M<C�IK��9�����t��]3Ԯ�'J�TB�*7�c���*g�7j�BB䉷[6�����?ꌕN�(zxB����a�1N6��ap�r�vB�ɺ`[n�AG�p�r)
�dݴϴC�	u� �9������	2��Li�C�ɇ5� �����$S��	�oT�;� B�ɞa�X��iZ�ݰl�uC�Z$B�I*�� 3"Q4�V�IR��"cB�I����L�.C>E�V���! B�I�Svhݪ���.}�S�x]Q�"O�xv��v��C���V�>�"�"O�%�C�2Z��h5*����Ё"O�1�Ӄ,��g��7*ݨ2"O��S���X<T����\6o,�
�"OJ�*a���Q%�	���Aꕩ"O�͘!W<UHm��A?�`�"O�eC� �F9�}hvlS� qR"O�h����E�D!Sa�ѓy�6<�%"O����+L�R䚒o~N�H�"OH�̖�s& ����X��"O�����vվ]�P��&e��c�"O�$�e�M)}z�����W�l��8� "O�倀�I4��|ġ�/��Q"O,��ajK49�����K���"O� 
I*�HJ�eN�`�Ӏ�l����"ON���9�@�JQ�;lrtY"�"O,8��	 9~��#D��{M��@"OT�B��A(*I{vC�C���"O�8j���gTj��0�O�<�{A�'���'"��'�b^>���͟8�I;Y�LcUb���9���,"P(��	�L�I��l�I۟$�	Ɵ`��쟀��2q���dlU�.�(�BF�;0T�����p����	��h�	џd�	����I4xz>��#���w�6�Y,�j�"%�Iߟl�Iޟd�����I˟�����ɜ,AxX逆�1ߖ�)r+7��IʟT�	ğd���������t����,�ɉ �()<-��ٓA�1W�<�	ǟ���؟X�	�d������	����O��p��!x��f���T�~��	����	ޟ������I���	�����<F
�%0pE�c�,L�bh؁2z,��ş�	�����L�Iӟ�	�� ��8iۖI����3����������Ip�Iٟ ���`�IΟ,�	۟���5#�z���B[R�iK�=�n$�	؟x��ܟ���ß��I����I�����g��M��J\1s."���?Rbu�	˟��Iӟ���������� ����\���U�8u�%gm��i�`0{#Hi���d�Iߟ�I����ԟ����@�	3L\6)�d�	a� �:��L0b��I͟�����L�	Ο����x0!�Z���ɽt�$�G���<(0�"B�C�"���a� ��$�<�I>5bZs�@d��'�����뢥Fx.�c�-w~2�j���$�Ac1��$�O0t�t$L&a��2����j�"q�O�d�4Gȇ|����BL�$��O�5�u���tqEƲ�y��"����cE�D�A0��5�?ѝ'8���C@&-�y��!Qe�ӍK3����f�;rJ�Z���-�hu&����'����������]5e�0�R�c�40�"�a�9~xFT�I���@�e�+�?���@�F�D�A�H �_w� '�٧[�|@�5!��X X�r��:�Dƾ^�́��(���[&_�L̓׾�8���nP�Yg�[��0T�󍏃a	�p���d/�d��(��8��$��O�qÉ �^\*����O0�dޣz������d�O��D�%<����	� �N	�F2,�X ���'_���+���1+��Φc6G�yD&�j�b�|:3��ܟqR�� n���p��
;OO���dJ��$0��#Z�8��%-Cܕ���4�s���'r�J�MG0F�L<���ӚmL���'�,�BGN�&������]�	$,�<c>YS��T)JE\�E��tj,�ᯏ�fj8�PuF�ꟴ�QFL*Mk��;AƅY�'!�7m���u�d�K��� a�l(,reC���]����_yBG�O��I���)%m
���O����lq�D�ԥE�0ZrE�2�����	�n� ˓���@���?���?����R�̧�?ɤ�4[�ѩ@��HJ7e%V���?���A���	s�(�c�"2E���2'~�(Q�h`8����j�`��s���f�>d�o]�1/h��Gf9r�'3�����I����򨉩~�$���N: �ɒ�OJ����O���O��į<YP���,��9i��h1�"�M#۠���	�O=��̓`���'��Y)�O��'1��O&�����;U[v����/�����ǌ!��m�ňR*M���-�̸�#w�1��c�'~�3߿C��J�l���F�|��`�W�j�*�4��?1���?���i�F�qL~�;#x��r���Wg�H:��T�:�n����?)��42�8z�8���ڦ����t1N�I!e�!�4j^�E|!p�ªv)n7�L?y�L<ON-�Ӻ+�����uwJH�*"���,D��(G]I�m��W!X���Ä�?�oW�v�I(�?�H�E$��`��ȟQD�>��b��M�?�(�����֟�IlybO[�O��U�'���'��,,N�q��&�/	J<�f��#N�|~r�>����?	���^?�#Ƒ�?'��S;IH܉��Cn1( s��r�~�1w�7��hm��2���?m�u��(Є^OyBB�SA���D�E%�6e`���,�D��-��� с�O��4�����O�˓Mx�����Bll�i�N�f�B�`�"pͺ�8��?IT�i��р���v}��'3xe�l�9xY��,H��ay1�'�v����l�p �� Z��y��UzU���y E%��<�A�->#����J7Q\�A�@Hӟ$��z�Vx���-�?Y���?q��u
��S)����h��
�  �m�m��9��X�7���	!�<Q��BV�T�|J��WC��w�H�ro���V�W M�e�`�'�bk ��~���0�0��O�N��İ�~�"oɍy�zŲ��M&?��2g��{���	��"]��=OjH��<qc�'~T��1!E�$(��k!�Y��j�
�ឋ ���'�R�'%�ɝj����S��ݟ�����0{��?H�|���-J�L9�'(�����+?2_�@�����Td���OI��@�ϹcHi�ԃ�14�8z�9O�hx0F�5L�7m�<w��'Nάm�fɖ���FY2aW�M �Dw�F,H%'_\2�'�"Ƈ�dV��Ւ�d�'Q�wy��K���+(���n�.x�I�$�'h�㥾��'7�6��O��3r��� �:(i�͔*4�u�&m��5��
��؍jgƨ�x�`#s���@�@�<�P��;$i�ם�_�ؠ��Dўh��aJW#��6s��0D�D9��2�?	���l����?9�����*P\�HTh OA�� ���m�ʘ�,O�}�1%J�1_��d�O�����(4f�<�D���_��an_�qH�=��j��k)�I����VBx��	+��,[5�?�X��*6���[sKfBL�;�4~�b��K�g3�ɿ؎��'��0�cA�<��'�)����~��4�l�#P0 F텧P�r����'��'���'��iy0w�O����Ip�D7�@:g���	 �׭j �������� V0�-���ʟ��I�<�X�C� �f<�B��Ru�L�RK$h4�Xq	µng2�r�LP����B�A��ө��� �}��]�)�x�8�CSa��Xz܉����O����O�����䒟�ט9��	���6)F	En�:Sr�$�O����`L �A6�����Ŧ���'c�d��"hD��j��O�h�ap%��=�:$��/����CӅH ��4�b1��o݉��F�<I��n���%�ZF��qi��n�#�&�O��:"f�ny� �O6�:p�Ȁn0�D�O0�(^X����%ZR����s���D�O:�Z#������?����?����&�@�h�[�T�tnQF��uy��y~M�>y��?�U��S?A�.M�j�S*r.� �:���#���$x���e�B�a���#*�";�"������'��-"3�<��nP5||BH��o"Ȓ��{��Ð�L �:��'��O��' 剩W�<�"�#H�#r:��ʇ�ov�����ѷt{ ���۟�޴�?�'Ft~"�>���<� ��"9=�:�Qc^�ѱ�'���]]�2��p	���y"�׽@}xt��L�4,ʖ�t��B�%̾9���ӕ	M�Aܤ�z�L�O<��	����#dL�埰������*��ŖO����'AB�:|Ё5@�.0��˙/i�xr��'��'��4.����'~�6=�PH��aJ�<fL{vhAN($ؤ	�O&�dǴt���61|p�ɟ^���f��b�Z�H-���� �����A8�.U��v�z�*l�(� +Cy���O����� `��$_J`a��bF�Z
<�2���{'����O4�D�O~˓f4�$� �F��?����?AՀ)$�20/
�R�U�UuF H��E��Q�'����?���$8��Wm+�T��d�����(�&�H󧫄�<ك̄;-@��ش'��`�,�"X�0:O�Z�(	��LDcW�Z�g���4�ө3���������	����ㅞl�������X��eT�VҌ�٦D�6{�t8dP矸	�.Ɔp��|�I��`��4�?���B~�w��K���f�Xm��@�&�S) �fl�Bq�O|�8�D�u�N1R�ğ#(�E^w^�A�U掜5�NX2��'��4��{Čܔ'a^�I���@�i�O"���OV��[w�F�R��	�=ntZ"��;x��o�<��,Tf����?)����ĭI�|���+.���oǪ@@tjb�H?m��q�0R�\�IßH3�e���Pb,T�����:��5k�j͗Pp����ܽ?C�H� )T���zA���<�G�M�"�I�d��'R:�$N�e(��4D���.�i�@�	��M����OZ���O(��<!-�(A��!�����E���� lb��0�L���̘��-����'d,}�O*��'���'bM��� n�Pt�@`7 �!Ä�`7Ġ��\�4�K�'M�������#7�Q�D��'��k��?�pU�!�1? �bf�*j>�1J�� h��'D��O���F���wN��8� )h��*X
t�쳣�'�B�'�ڑk�!-��D�'gr7��O �1�:O�E02�ȼK�P��L��}��l
Ç[�J"�$Z� ���c������\���%[�$�	7sF�Q0+Ÿ0��J�̵1ʕ$}�� ���Z�!b\��2�� xV%��?����?��H��D1���ÍZ�v��IY�?����$/n����g�Oz�$�O<��V�x۶�T�@�p�3%���s�9e��ؑ�OH�d�O1��O��#�cݦ��4��7�"\�N��Y�BP���Å�n�㰄��ƤPp'�_/�y��q@�����J��)O8�q�nL!V`�l!T��.��T��B�ʟD�v&��Q����ڟ�˟l�	By�B�1oj�����K�O $p���6����@(E>��'mZ7-�O��A���� �O^��!B�+s�\=`�I���A;���$E9n���R�6sYd���8OP4CJ�u���3��ΓrB�@*�� � �6�0���s�~E�ɛ�?�uD��#&�����?�����C˓��)��+���'�=C���Ȧ��\H��3���*z�����OR�$�BL��8���d�Φ��o$�E2sKɦ\(q�CH
2-fj��IğdZPi��(���K�cp��+"����	�~�a��^�&���ʃ��-lx���ʨ�y��>C�b(�V���c.O�p��Y&�"���86��77~ @ �K�0�*A�'�˟���Ο���Ny�KȄM�l-�a�'9�'����F��?:$�(��d�/a��d�'k�U�O^��'B�'@F�h�'a�q�e˸�$`­�0�@��BN�d1̓&y2�6���(`�1�^j��C���?�%�@�^ФE��!�0)�p����@;2H� ��O����ON�B�@p����$�O���Lqf����&on�;uhO> ;����4��Q�1��O��dצQ��-�v�Ӽ�3i��?z�P����dX�I4/Ӥ:�l���I+�?	�%ϥw���Zw���١0O���r��<�uߴ;;H%�%��e \H%hL5w�`I��	�����B��;�D��	ş��	�?u ��/Cz�R�e�^>]��Qy�%�'C 5��k��'���O�h�k�O��dO�+��A��G��d��+��u�꓆?Y��]��3����!BR��."bSd��1�Ā�'�Ͻ���C޴b��ʘ'���@�"��<1gM������ʟ\󳎞Q��d��^�0�^(`�fpU��ݟ`�I̟,��ǟ|�'x���g�.	r��'=�`� �˾]w�h�����b�w�r��w1��O0��'���'�.DȒ�\8~;�i�G�y[F�h��ߐ�{e�V��*ٙ�'<��`�\����
ћt��'s-7&���0U�D$�q�"�.���`���a,��'��O���˦���w!�8 @���2�s�,�	2 �'���'~����R����'�(6��O|u�a2O�P�'p� Y%�	���#%@�39���㰙�����ޗE�Ύ�]���|j�݉1
�5p'C�F�paDȅ��`	�b˓hx�̥>F|����'y"�'���[�C�)`�{mO�$�z��b�'2T�h�䒌�.�Iџt�	�?m��05�h�
�:��K�d�z�R)�I� �ɉ6���ɴz<e��5���;0��.x@X,��Q}��2�ᘗ.#Ȁ��`��+�8��;O��m���?��+�<3Y��8A����E�T}NH�!Q
�B���3���!���?!��|����?�)Or�Y$J�2����9[�|Q��U��kG��<ٗ�i�B���E}B�'RLD�+v�Y�$E
Z��Ͱ$�O��
 �U�?�PH���V�<��%(�&�ݵ�m��7O� ���v�Y*"�@#�&
�"�V�h��'���1K��l`�H�O��$�O��)��~�';0-;���3 xl�����8���H'��(��?Q���Ń@�|
��4���w`pC�̍KxИ�a�[->���� �'4��&�~�#���O�
:��`���+*�r�����	2�f��ˊ'd�Ɏa���0�'�.���K�<�0�'��ir5Q�V���0�j��7>��P�C�
�����kb"T� ��B��4��ѕ'R�
 ��1J�:����f�Q��2�y"�'����?Q�uE0t�N��L��B��@98��eM�0+R��
<S�@ �I�|���z&A�Q��y�f�a������Y�	�9�Du3�GE�JUiC��+(_y:4h�D��'|�!ޏ1��i�Õ���'���'eL�S�O�).�ܰe��Y\��0��'�L2U+M�1T��'+V6M�O� �w����	s"Ģ�II�.)��!�B�H�%�*gHv��� ��B�b��@�$�<)�N/1@ם;i��r�,��t�s���W*|�����@�	��?�၄�
h�0���?����z@�W�9��a�
��g?�\���'�XM�(OM��.A�.M����O ����d��?!��#�a��x��G�A�pHk������O����y�D�/C�8�͟eh��[�r:�����Y�0�Jۦ�[�*6�6��*lY\�	�j��9�5O8��@�<Ѡ�'Y�\��D� �}bw�	�a�HYxA�]�[3"`�e�'�R�'���'7�	3D�RHauo[ß�c��6ߊ]�3�פh���U�A��`�ٴ�?A���~~b�>A���?�ǆ]�Qm�qQL[�0�F�r�)�9n�*�M�y�ةvhW�<��cP(Vl��]-�r�0�Z>y��Da����ƞ4-����Q�j�@W�_Ȑp��?����:�G������ T#b�� 1�0?�ވ[ ���?���?���; <p�'�?Q�i7B����y��ʿd��X��%X��,�cG	�M�6�O����[F����,y���x�Y
/��<�#,Y2L�ޜ��Jل!Nquឝk�BءTI�O��Q ��Ky�H�OZm�vbA)Mw�D�Ox�D��j���g�9� U�PE,0�����O�ʓ���Շ�!�?����?��'�܄P��Z:�(��sB�+��)�o�A~2C�>��?1)�k?�QI��>�0>!�� �	\�?��q��Ni�L K�gK����5���Ry���T�WP�C�;3U�˓-����bi�"H�i��'�j��D���'|P�&�D��y����d�'HU�����Sf)��C�/���Y13Y�[��ٔ�����	��MC��H�4	�'Z�꓈?itI۬#|d�!4k��t�$����?y§˛m֦� �ϗ&����'8ҼY$�t��U��qM���H��y��G/^p�؃W�W�R�'�O<�{�M��ZP8��O������|��%t*,s�-�H�"tkے\pDr�	��?����?��'����'�?Q���y��w!ܥŬ	�%����n@Y�'Ě8c�'̆r�{�d �Q��;I�xț�L̵<5V��a�?���Ef�X�������dӚe`
ʓ(�b��;jzi���'�L ���[�`���'FҘD��'c��'!�\��`V�?
M�����	�z_�З �7"� ȕ�Q�!>��	�RT6�N�	؟x���\�B�	(i%��Pe��xIh���21�ܹ¢J!SH��W�+H�0��ϝ.p���V�arE��~��9{���1�i�6	��r1���g��P��ğ�B�J��q&?��I͟��# A�����I�HK"x�AʘX���).��M��L�����I��M�E[�]�y$�S,ԽQ���5V����f@r8�%b�,9�D��{�4�[w�=QA=O��b$��u����3�dP�R$D�l����ϺEw��rÞXy",�O`�2��E�A�����O�����(@�#��3A+65b�!^��x�N����\e�PU�O��?����?���ʹ�'�?�t!G�\� �˪V_�찖�N"k�I������\���r�b(���?� a�Ƅ5�����*_��K4lV����#V Ѽ�	�S��ahE�'5��8�N�<��'(R���+�2E��Ґ�Z3iP�30�Q�e��5AB�'���'���'��B{�����X1ƌ� G��q�NA�'��Z�S՟�i�4�?�'��y~B�>����~���L��t��m�<�\�9t�Z�<�B8!���+0���e*i� �.�M���J�/���j*��Q���Kdj�q!@�.Q��A�bW������=>��	ʟ��	�?���
	~�s�Y�%�+Xl�q)r L�eVp)%�ԟ��	ԟd87);{�'	H���'ndI�'6����C
�0`�������B�_�~��M}I>���|btl���u7i��Y��7BSܽ����obE+�,�(Ą�&+��yR�'P��I�?�ui��|pBr���?���-�4T���;S
����cơ'FL���?!,O��U�+w�$���O���韐tC&�x;�I5G�D�=v���qk.?aRU���	P?q��O`�������h�.���*�kW=?��TᄅZ�,�)�2� p�v����̄�y�'Q{J�I=,��.O�Ћ���e���@��
6C�u�J�|C�\�|P��������EyҫW�[F�$�p�
�7��"я�?_�j�gAM�/�R�'�B7�O�������c�Od��F�`H��I�:��r��?~��^&����� ��H9�0O�X�gb�b�i����3O~�yB^2Pl��5��;&Aҁ7�'�����,1��5!�@�O����OJ���8kz~˧!a��A�.���{�J��A�`Q�D��_�p`���?y��������|Z��f��wvx�燔Xt���eBZ@2e�'�§ع�~��Â|�B��O	��褵� �q�摒	rܭi���7G���,��Yd2扚.m$A{��'����Ӊ�<i�'V�  &B4uR��#�.�#UB�/������R7dC"�'3B�'L�ɪ��T�g`��,�	ҟt�Biê,�[Fe��Q�|�c�şD���)?IT�D�	��5�����q���D��rI�"F���0�̜/k��� �?O��h��t�H7�T�a���':��ϓYH*�3-=%�Tya�ׁ-��M�lD��'r�DG�w���t����'�B�'<�M�f"�@^ZP��I�l���`u�'k�A���I����'r�7��Ob$�������pC���7��ѡ쁏w��1z���._�����0��������y2�N01�e����� l�K�?R�D�V��E�Ha�:P���?y���[L��s��?���R��܀d�>486%�1K��$�2��,�X�.O��c��Oض���O��D򟒝��9���d	�T�%�&*]�z2�=��E̚H�
D�'���'j�,�'3a����J��Шk���S�h�jɲqO�21尽lZb��ϓY���
6�|��)&L�Ky"��O5�#n[�&qs��U�}�Ӄ;g���
���O���O��d�OX�3�y:�G��?Y��^�'=
(�/�+p��B`��<i �i�2f���dHO}2�'(�n=p��1� l�r�P�qe���^;U�E�������y�LT��%�;xs��2��|
��w�]�a'ȝ�x�B�ރ%��x� ԂvwBL6�'x��'����\	3���y��^�P$����*�<852�aȇw,r�'�b�J�irϟ�mZӟdk��p�|2Ӭ��m�d���3G.�-s�*M'3�$��hJ���g�O�4}S�ם�_{��ϓN�.�	[�i�PcUe�(��{�������
s���O�����M�����ڟ��Iٟ$��/1"�f��@��!W��Lz�/ҟ �IXy�mP0-��ԑ��'b��'��4A�*m:�8�Tg�\M�$�s��/� ��O�'���'}�@�'�X�ȵ���|ڗHe�kU��FT�б�B}7�A�2�l�+Cө#����#��'��2��ԩ&f�+iu��R�/jx�u���?郋=t:��?ͧ�?����1���&��Dp��ʄ�"H�����N�/;����O�n���$�0?!�X�,�I�N���M��
(�yBlп66T����	\J�Ռ �&�]�t,|��ġ�,
,�i����>OD��R���)��v@X����9$�'j���dT�0��"���'�R�O؊Y��]>-ZQ�����,��G�*�陰��p��ɟ��I�(�S�|�2��'ʐ6=�J)af��CSĸ@qe��Y>��t��O���L��dV�sU�*ȟ��3d�j��9w��K�E��B�[�LhQ�`%B�8]ϓnP��;e/�O�hf��Zyr@�O�Ÿǎ٠�l������j�-Z���"� <F6���O����O�ʓKlH�3�����7��O.�Dݕog�m{נ�/'���#�@��4���d��z;�	��d�O��d�<x��$�'(�9��(0�m�v�S*��J�Bۊ�y"#�k�`8ܮ +��(�Rx8��'���q�Ҙ�Qv�װ-b]j2
Ќ{	��I矄���.��D��J�������ٟ8�⃚�G�H胂A��FV.u�w��ПpB(&��y��� �ڴ�?���A~�wH��;`��,J]L�'��ZAA��X	|�� ��'@0�����j�.'(?�扐1�B�{u���S�hɀ�w�?�T$ҤJA3[�����<���'"�;G�^����'���Oۖ����S��rr�K3�!�7a�+�+�ڭ�&fZğ ��ן��S'orM�'?�R�Aƙj�ƨh�DI�yמ$	��>1��?���z?�%m�s#|�'W2 Bc,�"�F�H��1Y�`aG��1Ɩ ����<��	z��$�9��$�'�����0&z�eH�w������T���j�k�=j�D�Ov�D�O����<���(}����{�}�b�O[F�gnT���}�������'>��Q�O���'~��'��Y��ɓ3Jp��G����P'FHD�܉��Q�d�� [�'t���	Ӻoڱ1�ԁ�Oo���6�~�iu����d��@�.H�E�FP|�[�O�OT���O����R���N5���`&ؑO�n����AhS��D�O��D�oԆp�M�<y��i��� ��y䐵[��h@Ф��B0R@��ב DQ��'GZ����ڷ�?ͧ%�~HXw��1�:O��0t�U@zq�q�N��X�$R�p�(�b�f^�����H)�ˈ��?���?��i�Ƹ���"&B@3(��?����$�+IZ�؃G��On���O��)�b�`���24�@7�O���Y3s��P�O����8��',v`2���|"kb�($!�<3x%I��b>��Q�TeX�����<�ӣQ�@�$��z��'pZ�B���bS|P�E*���L�j�O~�S"�kC,���O���O|���<!#�
c!"$���	B��h��.E�rS(A�?1�T����'3l��O�A�'�B��bF�#b��8'Ǝ�q��H�L���
�8̱t*��Y͘�̓1%,�`��|ݝb���n�d*�~�rJ]D��TJJ�2M���O�,y�
�8���O*�$���4��l�|�b/�:o�Lm���R�>n�H�䣙ھi� 8�?���?���&�x��'�?�6��y�;{�VP��H1P	0giZ�^��'2���'��Bb��X�$C��_��n�5Nch��2JS&B=�*�Dq0���t�0X�&�a���W{�F�C@r��(wL�Q)��'5�I���zi�|ʳ#S� f�̺��'�b�'}�R�܋wNт	9,��	ʟ��	�N�8"�K�F,2(��_��-��e�|��� �	~>*��I�h�l�/�T����(���Vk��dU�z`~AzW�h�� ��|��*��<��B ^i~e�C㒌a*��O�='�\P��'n"�'���C&N]3�OOr�'lBm���D�#��\�
�4@��E f�"��v�U ��'y��u�|���r;�i�E��`P�y��
UeG"[t20�BE�i�P1)�O����ˋ�v����R���S�'��$�2 ���W��.S��`���,Ow���	�+r4z�B"ο<�'�Q���g��'�2�O�L���+�F�b���$Ds:�*�-��j��9`��̟�������֝�M�Z�S�����F����lO,Ď�`�������O��D�l��D�	S ��͟&���N�j*�d�Q�n[b���X%q�F6M�S��	΂-�>OB����<��'�t�aE«��as�7/&X�q�D�Pr(��A�'rr�'�b�'�剟+J͡A��ԟp�nE�G�8����h�x#!Ԅ:�����ঙ�ɘp�`�	���������Бsc��<	1Q��O��`2LX�%�&&��dm�ę9[w�L*��Z��G����*lU�2�.�b��,@<���L"N:TY�Ti�OB���O���VL�p���Q+4��A	��<}���2 ���O8�$
^mJ�a0�6������I�Nrf�ɒ"�΄�e��6�����I6}^b%)"����P@ț1P�2�4�bͺG�yݑa�΅�<Q2�Y�? �!��B87~�ɃS��q�\�9[�yr�T8v��ɰ�?�r�ȧS'(!k���?��S��跏��1�~����=VN]y��?q)O��qGN��R���D�O�����%��H��L�0&��t�^xz��,��I�����O��Ā ���$��eЛO!�|�/D�vM�$�t"�20��R4B�U���!Ȱ3P��ٟ�G���$��׮����>m�tgZ�L����N�� ���8�8�e���i>5�I�\�'rܘ�E��0x�۴	�Ė�0bh@�,`��P�2ڴ�?QS�s~�l�>Q�w�ظ5z��p��FH�a�mp��r ��*�mL��p���<9���.p��֝�5�戹�6Ox��G	Uh��`�Ŋ)aR<EA�'�����>}��҇�O����OB���:A!�˧)O�PH��ǙC�as�N�%���0�Ӳ3b������?9���J����|Z����w��aa)9��X�",���(���'VBhI-�~�琫{YZt�OH���r��$��B���L�z\AD��7v��0��`�\	�IX�D�R�݊p��˓XRb��'*�
��'�0�Q�K�P�!D7�Y���'_��'{bR�X���%�
��Iȟ��	V��ɡ��$f6<+���O�b��ɉh ��?���ٟ�ɱ2���	0dj��au�P�<H݂V��3>Ҕ1㗵 ��T%l�raf�05�i�|�@S�<��J�r����F><�����\�%�� W�'���'��@A(����O�"�'�"��.(��&��<�@|)���I�%17�Ձ�[�0ߴ�?��C~�wMF��E�,�" �P�Y�	1�t���йl�))`�Ov�[�
��u׍�#󄘸�v��\w��Y��j��W���j��٣w�i{� �,���'p�$��c � �I�O��D�O����+�l5#d��CYf:�X�v鈳�<��Jܝ�����?�����I]q���0E�< �GZ�#O����.^�g� ��?y�q�<(��$���Y�@'�b��'y�MJ��Gx3Ơ�TiO	:t!��GݘaЬ)̓K؞�۰��O���gJGy���O<�e���	��IQ��'�$E�K�;��^��?I���?����?1.OLh`k>f[��/J���A4�	r��A��4?�N���ڦ��I:eN^�mf�Iʟ`�i�yBs��m�8E���>��a�4M�Q*��,��P��'Q�9�4BZ�;�&�HGD˧22�-U2�@�L>T�xe�"�G�C󾜻4#�SDB�'���O.�����wɒ���h]�:,	��M1����'���'���� K7I��	��M����J��\4���7텧9v�Rt��
��Q�ECy?a2�� �nP�i>�3 IU˺+5���y�k¯X��S1(��K��7�A������
���9�N���E��4�P��c��I�x�I8�� ���
�gN�"� m������̔'K�ɢ7�T-[�R�'Lr�OANԛ���"(_0��#͋U`�(��D6���Y}��'�r�~B���fQϧ	�lL��L�,m
�]a�Ǉ�j���
Ô9�+ܴw�|p�b���<�����dJ�(��0R���'�N��%]  ; �'��Ē�*�/g�������'�BZ�@��F�N;��99�8�!Gc~�!(��W����I��M��/�f��'�D��?	��ߓN�z�����gz$�ybKӟ�?��.�0T���q�Ɇ�QJ��ΓN4F�@�a�q�Q���*R~l�Ї�g��K��ַU���OZ�Y2�]�E(��$�O��$�V%�tO�|BD�D���,G�$v���nV�h���(6���O��	��VO��O��ozޕ���N�U�k�Q�>����V�Pџ��	�&"���DXᅗ?���+�ĺ�Nۙr��{������c�JȢ�'؄�҇I��<�c*N�����|DƩzJ8�	��h�c�;��l���P�N~���Iٟ �	��t�',���3(�4E���'w����c���0�s�Q�	��U!��$�`}�'����_?�l�/-���'��	W�t����
��S �z��`�J��..����N�W�tʧb]���I>{�R��&�Ԡg��S2�G�sp)ύ��'���ӈ$��H����4�'�r�'n��#Eht�1JD�!��RT�'u
X���ÈG��' �6M�O^�Rg���+J$(����ս/���ܯJ�ңT�M���ɹiIDL kV��*R��yb���(M�������tt�Q�
m����E#kfH��'ո�d�u����O$�$�O��I�w�\�Sn�z����lDo�,�2�e�<I�jH7�����?1�����E6���.ob.��N�̔M�U'۟&G���'���'�����'�x�å^�d�Ӡ1{
i���dL�F��/#�d��N��'֚8 U����h�w�������͟���j�B�n!�q	�J�z��v�',@*L��؟$��ɟ��	�\�'o���'+��9��h��-Q����
�"Q��,�2�n���$T�[-�I���$�O^���$I�� �K³r��P�Q	X>�(YBWr�����S���dI�%!:� \�M�����[��u��,B.3)<P�	��x��Q`B ?�����Z����I۟�S�K�x0'?�<�N����4qA��S.t} |�	����ɶ=V&��q�{>�I)�M���O���[� s�&��'�[�8�(Tz?q�$�+D�D��i>	�B�Lປ���yrK	a�8�W� �9�'lP:�`�y��۟Hp`����4���ƭ`dp�������=^����V_�xۄD"�̖}�ʝ�	Ο��'�ՙ�`�4=��'��O���`��* 栫D�GuQ'�̃��DCU}"�'a"b���~�G3�X��'���Iq�J�jf���S��5k���u;�ϕ�I��GV�<���g�牠+X�l�'eh����T'W�2��#!W��k'��Of�a�K�#����O�I�O2���<�7Q�o�M�g�Ȉ���2�I��=H:�a�N�?�?��2����'KDd��OVx�'+�fF�	��Hg%�8[0(`mL/b`Y�e"��e׬T"��(�'[!d[��ەKOh���	1O�!���[�K�z�s�AW�&[���Aӟd�w�O:V�ȅ��������?[��F��Ŝ�'�����Wc��G��<��0a�χ:�r�'|��O��r�X������C0��IL��d����k��!�I��Hh$���W�i��'
Gb��vH�,� �]���3A�d�[�%� HH�(u3O�����<�?Q�DG�I9�?!�d(�\1+��K���
Y�@��M����� ;���?���?�*O�1Rd��z:����O��da�S)�(D=���¡M�'W��a��'�����O2��'��'�س�'���!F�ܨYQT� ��+�P S �>�0i�s���*b���Ec@�e
��?����s_����ɂ5|��Вqhī2|�Txu��O��d�O�ڕ��?}������O��$�	oGМP�
G�F)�Ƨۏ���d�k�"a����O���ʦ���8���Ӽc�	��)�hU�P�h4�40��X�qڜx��%ln�8 #"�ɺ3����yr)��/�����&��+��T;�R**���	� ̈D�X�'V�������7��O2�d�O��IUn��H���M�\�Z�땭��ȶ[Y�	9ft��"#ßh��؟��S-�8�'��Yk��Q/+q*�@탛$������>���?�t?��,�b~���9w�S*E�X�0DO-�d<X�!��E7(��b^�<� N�N�������'>��352�$��5�\��+�*�4بC��N/P���O^�d�O���<1w蔻@G9�����t��*D��R!�ĴDz���l��'O2AK�O.]�'/��'!0�$HQ [�5����[�.t�/٧l+\p��l��j�	�'�x|�fiQ�o!Fʕ�O&��zL�z/�4��%(�c��&�ry�TiK�8=����Ot�d��Ĝ��E-�9���Iދ4�x�����,^�x�t@�O���O|x�7C�/.���O�mZ͟��Kw���T��>:�i�� v_<l1�B�O�\�	)q.РSi�O�Șk�$�]�@M��pE���G�̕f|�Ѹ1���	�������}����X�<-�'����9m�n����O��d�O��S��%��`�0��,'g
=���OT��<a6&�/m���I��?�����v��4�i���'c����0����'���?I�?�m�X砸���h>Q3���(��ΖJ|bcbT5-O�M  L��RS|y�3�`��郆 ��Eʷ}�B�p�4� &�9X"�x���4���C�'Ģ=�t�tQ�����'"�V� �!�C�$��(�\%W�Z�k`�(l��dZbMy�
`�D�d�t�	���d�OD���.�żiXb	�8��QRN�O��8��^�;v�QQf� ��$�.;�a`]wp@8���	�<q6�a8	bE�;�.�Ă�֟�2�
�f��c#K��?!��?Y��+`2��.���'ψiĊ@�v��3L�d�#�A:-�����O|�d�O��I��|���O"Poz����T�4��0/�>�x�a��T�� ��ɷ^ԮrW�?9pr-�����&.	�5��H�?a��(����)��S�'��-�!���@A�"����D�韐2��M
?����� d�Y�3��F�����-?����ȟ<�	ҟ��'j��k!��}J�I�Ո�\���`�9rTq��*ٟ@"�k4?��W�@�Iɟ�#W����0��k&z!��.HZ��Sԉǻ0�,q�=O��"w!X2P���[� ��:h�J�$̵<*l�K6��`(�z���o��H�V�C�?���?ٰ*E{�z��O~"���?Q����h;�cD�)88���#�?s\�Z��D���N?��$�9�I���Ӽ+�#ߨ7�S Ăy�n���(��n�)r̆:�?�W����Zw�V	 =O�e ��"�u߀���H��u:��@CѰIV���^���d�͟T�患S���������	�?E�#�@�e>��3g��2���jޤ|�L�'�����i��	����Ӡ �|���D)��K�a�!�D 2ʱ�������O����4I�Dؼ �h}�ʟ\ӓb:C�~��'�V�r���F��Q^�7�+H[v��6�,�t:O>���<Ic�'!V\���M�X�ƭ�`��}x���"��5��;p�'c��'��'��I .�h\�`)����␶I�b�ڲ��6J+֙�v+j�|�ܴ�?Q��	i~m�>Q��~B
�]�`4�抑W�8�`G�VZ�w>J9�#�`���'�U\���l)�.������'*�E�R@�y�m{�Ĉf��P9�
4V������h���?�� &X_�sލ�5M��d1X�!(�;H�4蟴������G�X(���۟(�ٴ�?��(��<�*h�6��.9�~8Ж�J24��L��m�Fis-�֟�ӵ9��]�;	�H�'a~%A�!�=g�0�#mm7<4�h��� T?O`MCR��<9u�'�l��;W������ �I���q�L�hV*-E��)1���O����<Ae�e�lI
�?1���?!��^���&'<�rWl�;5b�eЅ�h~
�>	���?�# �m?��B�!�&�)s��s$d�<��ypΓ1S�ؔ��kQ�,M ��
Ȟv�j��� �'���a�N�<Y�	�X8$��4̀�����Gǌ��`K��H�AV�'O�O72�'��	5"�������;2Z��=�t,v�ZX� �������۴�?�`��b~2b�>�� #P�B4H��0�I�O��d����E�|P�@�Ńh�B���i��<Y���8�}�d��z��#�I�B+fM(��������E�O��ɩT����������D��:lݶ��O�8�hU���	�L�h���6�<���ƿgP]���'vB�'����0��T�'�&7=ﰹ�$�bv�1��RT�;q�O���qB�$��,h*5�ɟq�0aj�Ek��7@~�(��K����A�#	F�"�tOh���B�Ky�C�OTس�MK�^jl��� >�3�G�C�h�����MwL�$�O��D�O�p��հ�d��?��?ѧ�x�z��O�Vi�1��2�Ec�O�D�䙟��O�$�O�ж�O^�V Y	Ir,iR�Ŗ0~kܜ"�dځmF���'^��(
7�6j[�3�� M�X�I?I��4r'���0�o�>)r"8����?����?I�@D�!/���J~���?�;!��C��W*�Pu��&]1x�*t�@`q�[>����� aٴ�?�d�o~�w6�$ЃBɏYHmآ�ͤs��-fC�4E�d���'��PS¦ΔLM�2���,m�������`��*��t��F/_�b}� RW��-O���I  ;@Xi5`����	�\�ӛ��չv�B�]���q�f�DX��cu`�Ty�C��o0(!Z%�'P��'r���;��4�'�\-��BVD�Y%��a�,�)o�>���~�	���!�@Q>7a����� D�s$�6%->	�R�N�v�l�`�N�;��˕5O�0ئOK��?��~I�I�?�e%��Hj���ׯB<�T�Q��#g� {4d�?���?i���?!/O:M;�ͅ2c�*��͔,�����_�*ˢ�)������ަ��	)l��=v�	��i�q�0H�f8��RbM�L��p.�	�(U$//����'���Qq	ֺKg���˧j�7#@�k�,����_��;���Wt�rb�%���'�B�O�z������w��E�e�G�z%
�g\a����U�'Z��'1���(N�����'�`7��Ox,��1O~�sÏ�O�(dBe���f�ºi���K1����f���]�Sԩ�;�&���'�^`��CP@t!3��
R_X9�'m��3v$��	�G���8+O0����L������8�	e�V�{c�,��0B�
G	d��"<aC���T���A��?	����'�&o6p{X�D�1#a�,!�$(��*?ٱV�(�I�4(�f��05��\�ɞ;"+H �fG��|Ss��gM�a��Wb�Q!B����O�V�C���]R�_��֥�A�f s3�D�@o�:�?1d,ܵ?g��?ͧ�?����DQ�&�h�gfݦr�8l
�j/����O4�����O��n��L�p�,?��[����&!�8Dv�$��p�Z����I�Cnd�wfP|��H��v� �B��v��i��8p<OƅA�S T����"ǝ'(b`��'�:�d[��pT���O��D�O���C�o��'21H%��6zD�qO@�U5.�h��IV�9#���?9���2O��|���r8��wVX���o8x��D���8d�'��?�~�(��1ќ��O-�D�ֲ�B��~G�a��@�d0�M�&+�J�h�I�NJ*AF3O�x�ci�<Q�'}t����1�y�IÓvU�p-�v���rl�3�0<�r	��5�E���?�����
ǵI���0OH�u3�1p��Y�܈�'�|��?�����YyH
��L���磛^�P�c�E"Ga��� ~�}{v��M��֛��ID3g�D!BΘ�)5�ٺӔ�&���@��gl#��/wl��=O�̓��RRH��RՃD�>2��;�l�O�e0����@���O �o�����f4?ͻ4�X�AN�T��RCM�;�>(JS�-&ߴ�K�4�.�pA��?�u7.�s"�D͟f,��Xw�L�X��ȯd0���S̆u��@`��P!Y��'����Ǧ�4ۧ�4���S�fB3(��c�L�"��nᜐ"�O\��TB��4B��D�O0�����{?��4'�������AH���F���$�O���ܵ{��!J�N��ʟ�9@Nʅ@Ǝ%�Ǥ�E�5�ak�l��7M�L���I�uz���=O�-�*�<���'-^��f�#R��� HW�-tbE{%�B�G&"���'���'���'��	�N5@]��e�ڟ a�M\#}�r��ׁ�H�(�C��П8�ߴ�?����g~H�>���?����M���^�EA�5ʡ,�3C�l  �`��+���SN	&��8}�E�_w��dq6SW�t/��\����D"N�j�bO^�4))�შd�N��Մ�O��d�Op��M�MdF���n��S�Y s�@#o�ؔiW"�TV���?A�D�T�.(Χ�?I�i%�F��y�ąxzxٸ`�تF�a�W#�rL\r�'���7A���?ͧp�� _w�����4O����$L�Y� �j���b6(�q~H����"8YvS����T\��,C�?����?����-f��l�p@N|a�aR�jǡ�?1����dؠ=��6G�O���O��̑_�8�Dp��a��̜�0��h�Ŗ����O��$�O`0�V�On��fc����'���y*4�EvbU�Сؓ(l��'ń{�l�����y�� �TP�	V٢�c*O�J0 ʔf�S��ؿ;q�y���,��h�2M&������������wy��-R��>"D���/m3t�g�/1��	z�'<�v�f��N�v�������O�;b���F�]�vN�;~
�E��OHɠ�)�B�=��� .��p��Y�^w�*���I�<y�1p�$]Y`�B�v�cE ҟ� �D0b<+��W��?1��?��Q!�!�*�x�[ a/ik�Y���J�M$μ�1�N4v8$}�eo�O��d�Or��
�S�)�OR�mz�	!�A	��`�"�r)B�!H����	6���=s�PIr�?�땭ú;��&3aj�#V��79�����˅8h5���'�k$�
蟠cDc\���D��p�ƨK�4,�	�(4���;�Pf&�����	ǟ����'U�YcE�	��'eҩ��N����Ɉ>=aB��
�]�"AA����@V}"�'R�џ�~RbA�Aچ/B�-�V�	#��9�lE��)�<�B�}��U��׿SZ�a�O���ڔBвgϠ�8��U1�@q��2W ���W%��c�0�HL���Dr"51��R?����&��Ad�܀��݊�J #��Q�Ζ�]X�1��[��{�՝R+6���j��/H�0H�s��ɣ���X,���
��W����3t�6�(@EZ�8y�M�g�i�G��tt�� ̏)?b� Pw�ʴ H�=�H�t�h��v/K�� {2���r ��	Uc�3�m�)	#X�Y䆏E����w-�)�'�@�`j(��i��&ݥ[4B�P�̓�?����r?�s�is� V�i�%x�iTL> )q��>���S��䓝?i���?�ɟ�P+�c��.����7nӅjoԬk���%���su�ϓ�?�v��A?��۟p���4,lU8&E89�ꀱD�8���%�Uǟ<�'���'*�X�iw
�}:� Kx^ԡY�+ӺZ�F�iUe��qi�Ô��`�ɠ�B����$�O�k�b�OX��%!D�V\`1�G�L<�\��	a}��'y��'��	�p��T����D��^]�X��ś4���m[���l�\��V`��DG�t���'���U���.���q��m˰Q0�
<vj�6�'+�]���g�3����O��������D�BL�-�`�2P!K�^���G/u�'N���G�D�ͼ�a��
.�̹�v@Qfl�|R%(�Ŧ��'=��S�s��D�O��D�:|�'/�x� �.y�Ԍ�fk�P�6�A���>R�'I0T���&\��'ϲ��B)U� �ڥ"D��^���4w	�8�ıi�R�'���O^>�H�h�R� �ݙ���1��i��	đ`'�Hk&�i���yD���K�1���ą_��c��͑�zV�6���m�꟨���$����%���)I��Oh��ikL�A��O6m~H`D]�-j�ᙊ}��J{�'"��'=��6$�B�x���LWrG	�+S��6��OZ����SC}�i�y��'�`����b(�}z!+��ܻ��Mfn��'kt�8�|��'pB�'��I	 �&q��CPY:�E�i�,�B���ďS��D�O�C�O��'K��Q�b���+�q�7
�W�ܠ�|"�'���'��	�q~�4@�O�t�����(Wَ��3$�70G�t��5<&���ʟt�����'��)�O��a���bȡ �5?��s���X}�'���'��	���}�J|z���9/���ʀ䒩KR&x�i+:O���'����'�Ht�+O�i�O��T?��EPr�F-��l��x)���g����O�˓�蔠����'�\cF�IA���a��1��cxh�AD����I�(�<	s������O�s���@<��+�ZvN��da��
r6-�<q�c�m��"�~�����1Y��s���!�8��⃓�>�R*7���dF�ʓO���+��?��yʟ���W��飗�\�e�e[s&�MSVaB��?)���?����B-O���$5�P���,X�'��3Ee�
����Ο��*U�,��b>�	�C$ʼ��@�(�̣��Ƥ<&	�ܴ�?����?��@�5���!0��O�� ��i����
̂e�����я|
M�޴�?QH>�w]?�?i�'I1��L3��ߋ<P2$���M���k��r)OJ\Ju3���I:���O�X�JA č �"t��lS������>��w��I����	��X�'��-6�G]~�vnO%&m°e �?\+��8r���џ�xab����yZw�,*v#�`2>���ĝ4]�0a1ٴ�?�H>������O$u(�?1�3H� t���c��X�I�B�b�2����O牟o���O�bX>�P7Cq�.��,c���Y eJ��4�Ѷ�xr�'?��ן$�u-�B��'PT����
?�z���[����rӲ�I:s,����!��]>��P)�d�0ǲ��GK);ߖ�)W��P���'��	��4���X���'���5(��:	J���AÒys���6�R;H,��ɷb$��Dg����v��iExZwJ��� OI:e}.�@�ȶf���"�O��$+L�8�D�O����O����<	��^,�"ZЧ�ug��
�k�!tH����y��ZoA�MExJ|&n�� l�W1 PDi*Hۦ[d�#�M#���?)���:ST�X�5�P�H�'J}�` `�	F�kc��� �ΦM����ǟt����$�'1�3?�0��g���&�I�o���j��KN}���'���'����@ǯ<�2Aq>��1�7�"w�(���ljF�ˇt���'d�'���<I��?��"wT�Y�ɀ��3<�����䐱����'�L3)�<���o>A�ɤ`�\�"J-#���b��±��Hb��V�xb�'"���l�	ԟ��'K���7��A�p�7PJ2��0�{��ʓ�`8�����ʡ�o���'��	^6��@《	=ℼj�h�4k5�&�'E�ӟL�	���A"6�IO w�tAHc��ոeXB恢�@C��?1�$�ȴ��?������'�1
WA
�Qԍ��C�)p �A��>���?�����$Znꪥ%>E��+�'O5l�)��/I%ѦbI"�M���=$@���'00T@���	�O��T?���U���pF��9pf�MP�q�X���<9��c(�,�<�$�O����v��#)��v��,�7Ǜ3���;C&RE?Qch��\̓�u稍?�O뮛$8�=�%ꛔo�D�����p���,aVo�ʟ���ڟ����?��'p>)�R�ވk���!�M5�Z����J-j�B8O���CEʴ�O�OӸ�Hgᏼs%�ɻ�aQ1���۴̸,��?���?Y�'��U��IE�s=�P�#ᗘ䤸���RF�8]�I�N�t2��)�S� ��K
:�xp�t�2y.$�dJ<�M���?Q��)��JPU�pK�@w�����{�D7�\:5-ND�h(o!^�Ԋ��H>��|BC���yʟ����O�dMT0����A%N�DT�+�!}'��l��\�6����'oa���O����<O���Ɩ���E#Qd3��hh�
&\�h	��7?��?��?�)OJK��-u�Ĵ��J@<U2�xt��a����'
r��'o�e]�y��Oc��'�I��;��`Ybh$��!����'[R�'��S����z?��pC�쑥K a3@MR�j/$i;�i�:H��'gb��y�O$b�'` �K�'��i�A�ޥH�;!f�u�]Z��pӪ�$�O����Ox˓t��PV?�:��%#T���Ѳ�K͇� ��jq���9&��^�Z��O
e:�ޟ��O���u��J�t�(F�7�V|2t�i���'D�I1��D!������O��)�	`�L��+"�9�҈J6 X,PkQ4O�b$��O��D�����'��I��y7�^�f%�,@AnLF�7l���M#)O^�
sF�����˟(�I�?)�OH@[W��w1d%��Px�}C�MX��d�O�xb�I�,}:Oe��C��� M�oR(u�i�>`��x�^���OF����,�'�8�˟'�p�A�N��I��$��HrBp�#�y�a#��̕'��k����'�u"`� qi�\q&�R3cd�qa��aӐ�$�O��D��2�=lZҟ\��	�����ɱ�d�]1	d��.�7*m�1F�1My�7M�O��,�l��S�D�'2�'d���jP�A���!!o�t��S@�|�H��ָS@n�ǟ�P�V�X��s��S�?7� 8���ǖ�Z(L�2�� 4� ��R^�H�nk���'�B�'��'^"��>1�������8;=�Ԋg,�6(:ր���4�d�,M��d�O�<1�h�9O��d5	���¦�`����mW9~��"��(�������ǟp�O���Ac�pӪ���
�%~���0�E��u��Ҧ�	�ҟ��I�!װ��I�?�	��(
t�c>ט3wcbij�o� Lu2KU��=r��?���?�(Ot ²��F��'bb% oE�p� 8{xY�́[�`6�O�Iz9O��� D�O"�$�<{���;}b��o �aP�٢q�J��r�O�M���?Q,Or�)Mw��'���O�E8`�H�Y�l%zg��(@�X������y�Ӽr��'����Oj˓E󮅾	�n��D��-L���È�=�&Q��K�đ��M;��?����S�H����|�h ������2��%xZU�I��8�v�q�@&��	я9�	��7�H���˚-%���#�)a������$7��O0�d�O��i\b}!��yR�Ɲ}\�* #�&r_0����ڜw�6-�=^���O���X��|���� u�e���bƗЪ�� Nb����OB���330D�'Jy�'����M��ዸ�XE��?������Y�'�Rꓰ�yʟ����O��ċ8,���U+�8��a��4~an���y�&��䖶_��D�O�d0b7Ol����� ѨP�n1Z��׸"�]SqX�x*P�x�<��ʟd�	�,��Cyb$�Z_ds���/\�6�م(N�6�ybv��>���S�<1�Z�vaΓ�J���?�cL�3�L��,�M�Y��%P<M����?���?!���?�)O|���ϟ�|�Ɗ�7UL��s��ʀ_9�d�Ӆ���c[>���O��B�1O����On�$�&_|�ܷrݔ(I�H#X��]�]�$X�yӖ���O����O��F}p`1AQ?�i�!���:7�����2k2VaJ��v�\�d�5{U�d�r�����O0�9:Ovʓm.���	�1*�Rl��~V ��i���'A�I_�l�L|����i�h.As��^<����b���4Q���+���I֟8���f�0&��Q�w#���6����m����.c��QYڴ��d �h�o������O|�ɞqyb"�J6J]���M�2������f2�<���?�����<YN>!�\�S�%{H�9��ʙYu��+0j��9vb6m�	ns�Ym؟���ܟx����T:w�qbX�A)*�-�d�J<�46�ͽ3���%�ί�1�$�dɯnN�|ِ(ϒa�^L�W��v(lZן���˟�
��܂�y��'}�A�ܴ{�l�[fM�0Q�0��Ddh	�d��b�Or@[���Sǟ$�	�ܠ�إ9����`�^3����	�;�M���H�T��R�Գ$1O����C��s�)P�I&'��1����Y��d��>�pʕ���?A���?�+O^�9��>}��@��94��9�b�[��'�T|;��?���o�d�'Sr�Rw2!��F�V&�i�u�E�?�~Q��'m�쟰��ӟ��'�p�w>��p�\�ש�?tJP[���Oā�V�'�B�[��~�'�?��"l��9�FI���g�Rݠ�T5"�ȱ�U� �	�����]y�Cu\����#cF�c�=���0��qQ�צ-��0�n�	X���D�O2���5O��'���Ȃ�	"/��14h��~Y����4�?������\_]�i%>y���?���+;IoYHBfǔ<d��g���gqZ�	�����?D��<�H>y�9�xySǈ�S̜����I�v8�+'�i��	��2aشk������Ӯ��D� @^�� �F�1}�]k�n(m�Ȑ���'o���
���|��'�P�k�f��Af.�q"�
7BD4�o�4G*���4�?���?q�'%��I
.�6��E<u�Hc5��9q���A�^S� oZ�8g��IS�	 :3�c>���
:�D-1���;I�֐@�韊,
��Sܴ�?q���?9r$�1��I�|]���O詠�i�Q�$L�-��h�&'
, ^\�}nڡ��'o��'�Rҝ_��)���F�<{!�Y���6��O��c�[y2�G�|�'��H��M���`m��XW��?Ell� LT[�I֟�'E��'rB�'���l�����h�\��Hcv����X�x�Ƭu���ɪ+x��>���O(�;u�Z�SB�50nպ{�ȡ�6��L-1O��d�O���OT�d n^��Z6|��(ȀE1tU�=[©Y��9lZ�Wg��	�t��#���i�OJ��P�;��i  ��+�TYj�O�3��4��O&�$�O����O�����oZ�l��%/��8r�$P&O9�tr��
���4�?�uƈ�y�Oe��O�qO&��U�Q�v���E�Q�¤��i�2�'4"�'�j����'��'�B�O�
��ChԜ������qبI# ��~����?ɞ'c�nF��֝e����U��J�1B�3(�t�M�����ZX��$?�h)���&s�0�r"��
�eKE$D�� �J�39�  #��2 1v�����
��cI¶rd�y����s;� �[;+�L�ˆ��84&aXv����ͪ��_�=4歘�CS6�����߳p�����ӑ#)EQ��_?2O�mk&�T�lV��SAV�%C2�<o�f�����V�o!�Pr` ֛I�t!ꒄN>	�ݙ�.G�n��'h��'W,\ t`A/�rG�MI@�!f(_
E�[�G�~G �w���R�j��xQx��=^W�i� ��:����%̕;|��䄐<��m�4�ʦG� e��ɹI)r :!'�?�T���!w/��	�8�����Od�=�-O�@P7��O~�rb��1Bq�\���'���I;�f4�`ύ�<��0��ʮqk�H('G4��?�̓��ď�n0�i�vAT��,��(��іa��z����O�d�O��b�l_��^��l>MT���:*�@�� $����I� x�p`�+�ox�Iuc��=KN�	�.pR��6�Z�8��i�X��&F"|��4�:lO҈���'�r�טg��wLՇi�\�{��@�ўTDBk
TKTh�@��)��PX򏛠��OE�$ �6s�ڴ���:DPB����y�B�y�Q����
	��Ο(�O�Z�[5M
4V�-Y�	S<a�L�)M�z���b�'�'?; �1Ê<&#\�2��O���# �-�U���:���8P� �)��������qIt���o���*eq�D,�I�7X���Ңg*�
����4�Q�P�M�O��$3��)@D��F�(+di�d�W_&�IX���%�8|,�xVm,>�Xk�'�>�U�~z2�Dh~�^2���)l�\l��H�y"��kq\]��'��Y>q�Č����� 1s��C�L��'�R�E�ƹQk����h"�ԡP�N�?��9�&���M4��I抜�w(���U�3�$��UG�-S&�;B�ͤ�"����"~�	�@�������TŢ�y�C%a�~3$���x�IR~J~�K>1@D�=(`�Wd,:��B��`�<EG�!C@�����(u0�/�X�	4�yr� ��O��:O@�����G �g��5Eԉ+�f�O$��Q�R��@e�Od���O8�<0I�����Ob��R�G�`^���E�����~�ɕ��>�����`w@!��.s�1��aSh?��Dx�x���f��asĞ�Pg�MK�%��,k���O����k�>$��N$ONq�TmL/7ab�c����&` ��I����pZ���GB���"<��`̓*�x� H���r�bv(�9�ty����Ue���?1���?)�J˰��2����!2-�X%P��M� 1��qIV���$�'�L���	��9�m����5Ox�]�L!��/�O���`�'	� �
7:����Z��Z�B�!�y��5fA�I�	̐h燳��OXxD�$h�.F��0�e�7`�\0p�BH�y�ի��'��)��%źYS2�';�S
�~i���=v\��@�J��,���_�f�.i�	�d���@ e�j@�3}���?�p��pw�8%�͒=$��6&JS�'$|��çd��x��LZb	P�ys�Y=��<�3`Y��LD�4j#un:��g�� ��!�5 ���y���<�uH �߈S`�p��B��d�|�����3D��-#k����(V%z���ޟPF�ɷ��j	̟��	h��g��U1R�'��ʗ!wC���/Fk�h
r!G�p���/�0����I��	3�(�� @�L
)<�ȼ������܃B� �O?�d��G;�5@̊K|L�A�HB���d[��O�b�"~�	�Q���Ҋ��T���F��(&C�I*W�pm���V.|��ӓ���NO(�͓�^@Gx�'�yI1m�>a��.�,OB��t�	��y�M��r��4:7eS/'�AZ4��7�y���<Ko���cl��ƹ�3"��y"F�=L6$AR,Jzi����0�y�%� ,A`�A�*r!^H����y⋅�B�RMkS�c׸̙�V1�y��[�� $��<T�rT��yr�CP��l��K���i�a�R��y�#ߠ��ڱd~��I!6���yB  R�P�c���i��ͨ�BK�yB��~N��ǎ�[$<��נ�yr����8���	�F�:,�y�e?}�p(����$^�1āL�y�"�6qz*sR�I(2�<�i�H��yr'�\�"�h�+R�z8��䃐�yd�x46�h7�K&5����Ǔ�y�(Q��	�3�J
���`��y�i^+�=Y��^��y)��^/�y)L�Ԡ�)�S!0��XlD��y�\(��S�%�#���3E��y��/WJ8A��$ԋ��5��Ӳ�y�j��bQ8�dз�(��m�(�y��\�ȽBD�ŜI@I����y��Z,I7�Sħ�Q�p)��_��y�k�:���@lKi�<	r���y
� �)C��*tlP :XK��v"O�@��O#��Q��� �<v���"O����L��2,���e}�m�d"O���G�Z�xAz$��n�{�(�h�"OD���@��X�`��NG)�0&"O��#1��D����N�#����"Or�zqeݧ}#
�����)��	ڤ"O�!�� A��Mr����S��\�C"O�\C�i7C�DՑ0�S0��&"O��1f	�F�h�
�U����ƨv}������ը�@��C��2A�z�B�"O��R��N���@��a���c�x��f�|�'	T�c�mHd-�,`W�G)���	�'�x�p��5����f,Qv��xӊ�
cw���^!�]���S*Z�p�8IQ�z�Ǖ�/�'C�DX����ڇH��_�N��	�'UJ���EڬdS��B��E/*�"�`�{b��y��O�O�吇�G�kq�ɨ&�ݾn�	�'��`)�5G�4�i��[f�֍x3�/�ɸgQ>˓^xP�Q`+�5W����2d��,�ȓy[D�g�$`.����*G�Qϓ{�a����f���2qc-�MK(�y�@I�W���sbY!j�`����y�Å?=��q8w�f�⁻Rf���yRAA$>H�p�$ȆfG��R����y2��I��5A֠\=�1
��ٰ�y��*(h����Lҝg�f큦̏��y�I�n��R��X�X��A.��y���?���j�E�X)���2����y�G�$ E��4Kg�BB J�y�T.+`Yp'.B.94��Ɐ�2�yb� �x\�E�T!7���f�0�y��;��\04lB2;���(ƪ��yB��u��CajQ":�J�)�g	��y��
�!m��{��-+����E`җ�y���
�,4�)�:",h�%�C��p=	��8�I�8��m�P�z�	e!�x(�C��4 m��4�9Z�(
��Tx��x�EJ�S��+N���r���z\Ft ��W�ov�C�	�7F6aC3A�:F�&̫4/W��L0zgl#�I�P(L#|�' ��KяD7K:�R H��$�q�'z�i�U�ʟm >��]y	>�Y���&Ŭ��
�'��U;�k9\�
���	X���u��I���e ��E}�@L���bƖP%X��E��yH�L�,�2jӧ~�jq�1�N��'jp�5�^/x�#"� :_{��c!aʰ1f5CD��^�<� Q x�tL��e�Y�lb��;^���E�>�To#_��>�O��g-�jj���=d�^@	��>�!��V��<%?�2�
l�*ٰ�ʄ�7n��0���I��@�Ҧ�-{(L�x��'��UaD�[�[�n��clz�R��?�dhj��Oĺ�����U������	�y��F]rv	�Ƚ;d���eĘ�Px£��@�����	V6���hDm�)+�|H$�Z�[���� �T��z�iչO	T)���"��#LB�) h�b
*Pu�0I˓0[`��'������qEΑ��2q��:w��-Q��>dX�l�
�1���p�g̓|���q�.|�HX�s��HՈ0�ON���ѕ!���O�Oy,y`�Y��T�jff#,I׫�d��4��G��&�v����y��	92�*@��!��(�|��	�%��(̧.���a���"���Y�Q�,Z�M_R`h�IF�Y/���#;\O��#V�Jfy"Mީq�i�d��s���S���ZHf�Zw!���M�g�R�~��T�R9}��iP�V��D���R�]Ƈ�
'qO>�Bc�QG�S��rT��:�G�6:䤑d�� ��M"Cm�>��/�Gta�Ö�$/���8{��z"D��
����	m���gP�T(Јf�H� 哴J���q�M�<��4)g�����S�fJ���$�[�b��	<*B��	�S�H���T�w��C� 	X�R0zŊ�;*p�	@p����P�g��8�� �� A� �]*��T�\!��Q!�r<��aʇv�JT��(�.ʓ�f��C>=�`����J�4��<�y�6*� bT�T ��ͱS}f�A�21O�'rnZ5KS��%���#�	¾ޘa��I�v�X�>)�L�3,��d�c@(b3�� �rO$<�F@Z�y����!g��$>) �R�!&|��n{��V��/cx�@3�`[�I�x��O���� �)��V�}���jT+έ&|�P��˨B���]�Ļь�2
9�`�Jx�}q��F���O�|c�e�d��� �ۧ0J�w���-X�	+l+�!�a@$ ].<�ՊŘ��6-�;K�zM�b@_��:y�F�՜�b�����$��>� !�<��h��%��6�[��X��H�o��\�e��M�`��O��4x���$�,
B=`��0+�*�J�C��/t��X���*֎
�a�X��F�ݬ�L�S��<a��d�Hjl�d��8Xl�D�G�n0� ��-����x�l�#"�(�2a̶������ڟ��Ed� S��mY�'K��Э#*8���Ī��×��s���'	�!�㉋O�~5��I���%��l�1�đ4,�b��Y'jex��n]<	Cr���ODP�E��:x6���^�`d�Gx��"��:��L^��m���K]�	 P���2k���α fb��!�$��L�  1W�ө@CHyӱ��_f��ɰ23e:�0��]�\8�a��O�,:�fA�'��IQ�ρ&���d"O�(��&�h��[��Z�*`D,����"�?�¤P�!2�$�NԢ���	�{�,���iP�����q�����k���pGͳ-vv��eÀ�Hͦ	�U�-
�R��fo�,�����#�Tl�S��PF�S�)��^d���`G̞3�6�+BHc�(��������.Pİ��ޙP:�ѹ�"O((ɒ"�!!���6����v�'���S�J�.��Q�d�ɞ G�?� �'�p�
��'8@�E@W�X�<���ڬ�p�a�gsh]	��0I���9f`�r2�ƵP����HOҹ3�+~��X@���?�h��c�'HR6M�Z��YJ�BܸS�"꧌�!j���.��Px;"B�>J��d��f��X����c}& ���^$�nG�M"b	=O<H-ZքC8K�r8֧��:C�<��D>N@.�wDV8`Q>B�I&-�tT��ϴB)��¤��A�e�VEW��M)�j�O}��	�O����k�eP�₺U������.Z��2ͱ�	�6A��s��Y�mj�4�7m�O@h�%�k��آn^�>S�ͳ���,KRN�ÀJ�18�v���燫7���
uF����S�_.�Ɂ2Â�S��:���$�)�A� 5�������C9����Ot X-͎<#�M�%��I��'�剄;��	*�Ѣ(�v�EdZL���>)���w��6���c�B �!�L�\^%�V�� T޼�� �	'����ҋWJ��bѻ3�:��5��u�D�K�n,���n9�H* >D�Xx�.ٹG ��؀jL�:�\�5̋�Wmj��M(�5�G�еC��g�'�мZsJ�%ЮdĆB��A��[�D8��t/�9���L9iG�HjF��#�+˚#~)ȕ�r�'u��y�/\�q;r���△4����$K�`��]�� O�^cv�Xao����k�X��ȼk������=#czB�I�N:�谆ڞbʎ��oB�s�8T��S�N��+��X
 y&�;Ä#��<�E�@�݉Q�Ѧ�Na�a�J�<���(JO<��	E�*'z�s ���������PE�v�G2<�g�'�<#NR>~Ĝ`���@�\��^���Bץ4Ǟ� @��5�Zћ`"L<h���C�@��XX��%�O����M�5<4�#m��VF&)����%;� ���>�xi*�O�>-�'�VȘ7!��.�:�B�"��M�ȓ'L��0�TS��xBT�͔&�4�x�,ܐJ�H$31�%�MkV𧈟�ń�/�nTQ��<?�p����y��4�|�hRb��������$�֟�jVj�_��������M�l����9�6��K� �P����A�V�p%���u�����) .�t�4o�M9�}��Z(���	�J�*4s�۽9"4�$h1-�#=iE�G7���{Q��>M�
EP��?5�B/"[*���������;D���@ɵ��wE^� w�yPF��O�]�d�ʟ5���H�/�%!�ΣR�b�&E�ytL�#x'�Q�����y2��~L�[�&H1F|Y���(m��O<�hT�Uұ��'�9R�^�O�c�[�/"�\��'r��i�'��$���)s���
��� �%h�O :x�ѻc䏰,L>�˱"O�$Z��[a���IĂ�(.0��"O �p�e�3@�4}{q#G�=�d �"Ojj���h���!��x6d�s"O��b�aK�n�N���H"4"O�ݠ"K��(�;#P+uP��"O���������a֞\����"O�H"a�%t�Q�
�\n�v"OF�Z�ʀ;�����/߶A�"OX�!��+X�~�WM��d�Xi�"O2�@0�	�ifa�f�<�$"O
@��_����g��p'.��p"Ot0�f!�v��Qa0��&I6�|@q"O$�zU���"j*��e�+#�p�d"O��q�H{f���#Ϫd��%"O�i)�%J93��u��ۀF*$�6"Ov}`W�è%+jD��Z�(6��٠"O��I�$T?W!f�襏� oB8xk�"OΥ�3��BD��U���Dd0�"Oj��x��*a�@�XLj�"OR��P��e��
S��9w��˅"O}���F�o�d�a�ͯ�4�1�"OER��Y�+��
�B"p�H��"O�A�Eo�5�$=Y�,:4�F�"O$�C���d T
L�1w�)��"O|�:�X����qiK�w��Р "O�t�"���-᧩"	�>��0"O��ыK������O��d�R�RL�<��T�����F���S�YH�<�0��-F'���Fd�8u��@!ϋB�<i��1�HP�I�	f`ri�f�<�$�O6��D�"\>�3c)�c�<YA�2�*`sPO�
ht�Uo�[�<�ӆ�-]j�%ИS�A��YU�<�'&W�82�35�Z�k��RU�<��'[�]�ԕ� �ЉX��YYW��k�<�1�DP�u�A�&qT�A�d�<��Jزlˎ͉����2v�Ip�
d�<S�ČBV�d��LOr���/Vh�<�3f{R(=Y�PT�����Z\�<�2�٧@Ό*�֘N
���p �]�<�j�&"Z������D��9a�ȏX�<��6N�h���ːmupE�T'Eo�<�����~��qccM	~ҠD9� h�<Y�.�m�@�;rϘ�V�(�p��L�<)�;�F�A�N�$�����*�K�<	с��^�R�k]�1J��kO�<����8���Iƅ^�!s�`��k�S�<Qg
[�Z�<`���Ԉ<�,M2�MW�<�� V�b|��bOi��L�TEST�<QwH��|�.�SB�^8�xԙ��Iu�<�G�'b�d*1OF���({p�F�<Ia/[�J�43�<l�T�A�X�<��:9���F'�8R��h٤�T�<	F�}Ɣ��n�p�6�����R�<��kO�nVI���OBi�5o�N�<���Ŕl�ڹy�	�,n�b�ȑ�a�<��Yθ�z����8H�9���D�<����C�a�K��{�q
���V�<I%�rF)JnZ����ӡ�V�<�$�O����F.�$ A��\�<q^	�"%���Y�Y;ڡ�T��m!�D	B�R%�S�rQ��yu��<Oj!�\)�Q��M�>R'bD��\�4R!�� L�+�EZ0#�f���@ާ��`"Oq��O�=��H����0�,|AU"O���w�.]#��o��u"O�T��á��T�a،-ݴ�Qt"O��a$���G�.P�#��L���!"O`YsCO�� �3i���"t�!���RX�8b3��S�P��˜�w�!��ۨnX"�	6 G/EU�qH3JL�eo!�$�%I� 1�/X<7������0F{!��x"�xQfX�\�1�R1w!�D�,;V�3תnw�Yۆ��6E\!��-	��sq� G_r��3��
T!��*]8��u �=\�!J��B7XS!�D߲P���P�7P�{�Ε r�!�d�$���2 Я$��A`NA�4�!��V&]�p�1�C�hk�� ��S�6Ƒ�X�Ó.� �F#F�*G|�����r4��?�f�2q(�'(J� �U� 9c���	w<y��R�
�"\�p��ZѶ�pOD����<�t��y�łQQ�3p�)0��f�<I�۷R��c%�sZZY��al�<����q�H4JPƎ����ϙs�< %޷�V9Re����Xq#Nn�<��˂8:�u S쎮y�|��dm�<����+L���y�'7��(R͍l�<�׃�D��;�R"ܾ�3���A�<���[�>W�E��Ǒ�?���s�Az�<a �pJ����v4�T�JMx�<A��#���
�H��9�z�r�Nm�<��đ�#���Ʌ 4X�c1I�l�<���O�2ވz�8G�&Us�#P_�<1����2]zr���1G�
Y�v�U�<��d��vmbdK8]􂭒VMZ�<��!/2�f� .�<s��Ŋ�L�<Qf��_��h�<EX�V�KE�<�DD�����5s����aC{�<)@@�}`�h	�	+����%�l�<��Q�6d�{2l z
�Ѱ���b�<A5Bɮ2��}�R���P�8�L�X�<��w��P��(z��t�L�<Y�Y����hA¼[΄��t�Q�<���f�Hj�-9~�)X&K�K�<a���>�HH�5�O+>�R��ECF�<��KU1V��¤	�?��(]�Is�@!4�×u?Z
��7°jW`.D���K��^)x�`�+��)��O,D�0�BE]!Q-X�ڤ�9�N,+��,D��0���:)�$Tv��2OY$:��*D�tY#
) p� �K�vM��`��-��ȟ�4irbX�X7�k&�ǔ�b17"O�a�d��C��p�eԤV��UE"O8�ׄ޳y�Ʃ8r�K�S�.p�"O6��3�D�k�-
a��l �q��"O�  %%�FP"�B[�m���4"O�岠��(}:X�{�O�7�����"OP��T�,4��ժ������@�"O��3s�V@��X�'��9a���K�"OT����6
����E�ڥDŞ�	Q"O6,@�æ<��(��ڕI��-��"O�y���ۈs\T��"5��{�"O��'K��I�;�L)���:�"OB�P�Nݳ[�R��j�-&���H$"O�Ɂ���C��U��:x��4�g"O Q��9�,$ �'DnN<,�Q"O� NH�VD3yzl��Ft bآ"O�h�wD,�������.���R"O�(VǑ�ےc�DfԽ#a"O� {�JM0 ���ٖ��3`L���"OV	T�ׄLd�dKAtD��"OZ�)�/o�dUSs���"M�袡"O܀�s�;,M��A�.����"O�T
-G�S>%hr*�2򬬊"O�c��z���Ke�֥|�ݙv"Od=ࣇgA����)��|�u"O�9RiT�<�	6�v�n88�"O,a ϙ�7��{�jS"I����Q"O���	�z�1C���5�d�"O��8�Mދ7�h��؄�J)"C"O��г�˜5�	k$pT��["Op]qUfˆY6��'�B-���w"O
�[7���L0�P�e��i��p�"O>�3�D�O�h`Y���(�(s"O�HJB�A����3�Q	�H��U"Oh���
�=4| U�����h�D"O���q�#��!��Td���"O��@����Kr�(���X7+)DABb"O�%�cŞ�gu���Dی]<�0�"OF*��S4�̔y ��>#8�0T"O��cdS�55�,��,E/)�I���	[����65.�� A�1)�1a��@j�!�>�]��ς�OZUF��	/!���`����O
	�D��%�;b!�I���6�� �w���[��%�"Ol��� ÙJŊ��b�C��%8<O�#<Iތl�}	��ӳ]K�M�d�<Cn˘c�H8�N�9�F���nH�<�1�\�0cvI�C)Q��!�%SF�<#
 J�:��V�ۮr�8@Qu�k�<Y�*э0	���2�D�u�Ԁ0t[�<	 �3F*�\����c��0 ��D�<Y�
��1���X���<�B Go@x�<���9�t���O�qPplr��Z�<�~�Ndy�]1���ɔ�Z�<a�ǂD���ԭh�(X�S��T�<ѱ�Pxx�3�mہ:�)��O�<����7۪�R�_�Bz8�b�]H�<��/J�xQ�B�-���N�<)��-2���Z�Aë��4
p�Jd�<��w��#oX�Y���Yf�V�<���2�r$�e�E�ufl��P�<��N?{�|���I��qV֘���O�<AW/X r[�H�3	3PМ���J�<	���2&�@��D1J�r3��DF�<I�<d�&��1�1$D�4�$d@F�<	A/Ҷ0;���!"�,+���A�<a AԚ9�֤�&'�n�4�C��|�<�"C�B h�k:t@GG�t�<!�̒�BB� Q�܈97� ��C�q�<��j�:qՀQQ�b�BmA#+�C�<�(��U����c���|M�	3dUB�<�C�����Y�LFL��D��.�x�<�\�;+�ъ�I^�H�cZ�<��J2B� j�>09�=[���Y�<��G.@üɣ���W���R��U�<��F��D�K�N�IǆH#2H�<�ǀ5�
Y(���u1hl@o�<�PD�4r��(�`P�%~��R���g�<q!n��D+xn�XA��Jq��k�<� 448� �+LR<S*�;�f�"O�}'�H ���I� �@4Õ"O�i��+ί*q� !w�����'"O��r�����E� ���"4"O�EZ�)�;F�a	a$��yb�]�ƴi����*p�������"�y"mG)��Ci��e��Y�c���y���3��ˉ<O�.�#��y�DhIt���Fƶ{f~��*�y2�X -�.� ̇nEı��偾�y��.(q脫f��_�X�cb`�8�y�	��)��ę0kD
G��H#r�[�y���?�����@+F�X�q��ט�y¦[r��8`�VvW�)E�1�y�T:�6BS�W��!ed\�y�֍~�\��
KI�����>�y!��n)�oU��8�4��y�C�H�����R0]�D$���yRe��d����&��4i��ci��y"HH�_)N�R�+^�L��i�����yb�T�0w栀Er�����yb���\�*���K n�qt���yr(�n�쭻��>�jg`��y�DO��ĘR� ��ޱ��EO�y�K^�'�he��B֜s����k��y��)3y�u�$�g�j4�VaF�y�]����aiE7c�h��J_��y��֥o����ԛr�4�`iݵ�y��Cj�� r	��n8��7N���y�G�J�p&H�Qs�9��K��y�!d��f�R���Bl\ �yB�\�
�ȧ�0I}��˲�һ�y�Ă7ӄ	���D�k��i���^2�yB�O'w�~eXge��c�4-	D��yF��i�D�x�)�RV��p�����yb'�2*�a�����Ko�|	w�B��y��r�I6����*�����1�y�Ǆ
|����<����G4�y�����*��BG�y��9)�aH��y*]�|����7��Zd�l[7�y��H�p'l�7��U7*M���ۀ�y�l����CB�L�@)�����y�뜼M?:Dhs�إL�@)���4�y�h4���qM�D�v��p��y��W�1��u#�OJ�2��lJA(G��y��/[ ��n�2^Hq %��y��9Z0�Q��:]���R���y/�rX"��XKX��)Z:�y�#.���aDѹOr�#�߭�yҩN)T�<9J"��'���AmƳ�y�
�' ����οZI�9��g��y�چ(�|�e��~�b��P�̓�y�E��+��@D��)}Uz��VD�y���r��ހ*LF��gnӊ�y2��fP�P���;^����+�!�f*�B�ˋL�8��*�!�$�+�:�%����D�_�?�!�$��+X�X�b�٩
�zA:���r!���9M�~X��f�;�@�QO� m�!��
;�0��eB5ɒM��n�p�!�Dϵ���ڥ���6�Bb�TO!��l΢�Y&M��=� Q���a[!��	2(� !����d�P�勅�1;!��44ɞ�`�-� 	���1Q�R `#!�� ��wL�+4���2�Z�V�)C4"O�@�	�o^��n�NN��5"O&����;^a$�����@6$�"O�jQjN�S�YZ",�(d*�aY3"O������s��`@e��"�I �"O�I�P� q	vu�w"O�D� ��t���)M�n�Y�"O��HwlB�\,!e�5=�8Iӧ"OVU��X n���T�N�i�"OP����O��i��	RM�˅"O0��т��l�]c�- �,.�H��"OД*ګ8Q@�y���!-�h�Q`"O<�	���nƑ[��5M���"OJ�����d
��Ӄ�*�by��"O X�Be���H�@�A�/���`�"O�Uc���)F�0�fݽ�ưS$"O�eɖ�͌�Sr������E"O	�1�B�X5*��0���y�	\$t��p6�P�\�mҮ�yb����Ѕ��of�ˍ6�y��!x8@��b�$1��(� �y�ˡ[�B�Zь�%�L�uEۢ�y��^�`of(3�/��}�(�JE��3�yR�� ��x "�r�&|K� ��yr��
N�F��LU�{��ܫ�����ybn1S�&h%�O6y����u����y�n^�9��yS�H�mE�	5��y�Y�5Il��❙h|PqT���y���#}RZ���@�*6\& �s�I��y�
���CGG��p1��\��yb��Z��eх�����N��y�AQ|��4@�j�`���4�N��y�M�-���@��\ĵ�����y¨E�<Ƽ�sU)
������1�yrM^70`V�CrJJ�}�@$ˡ+Ϸ�y�� ��E"2�Zu�� SD�J/�yↈ�sP�B�f�7hA�le%��y�KV�\ߎ� ���!e��dQe��)�y�%�;"���l�[(&��F���y���'n���S$Xb3��y��r��a!�m��J̤M�r��	�y�قq�lC��H��Y����yb�������fg��=�:��G�Ø�y��Xm�F�SJҧ-j�Xai�:�yr(1B�=�"��6(�t9�!�y�)�8?�[p��5)?�0��nQ1�yb�֭[ذ���5LTE�w���y��!z1�UB �� �D�C����y�k�@�`� �U 1�`yG�S��y��Ld�B)��"{Il��M&�yr� 5��.�vr�lU�9�y"�	4�j��2�I�p�L�Z�O]��y"jM�R	�fz��:Չץ�y�9|E�]b�mڣYz�HpGJI%�y�-�L�0�i�C�M�lL�����y���dw��C�G�V�����'�y2	
~رh4e
�'�Tau�B0�yr�K���MУ�r�aQ���yr.X�0m���hԞ�c�:�ybE h2Υ{�FU�)S��y2C�/=�fř�jMst�2B,��y¢I�"~�{e�6J���0"ԋ�y2�ll�A�d�"A}~�:0)A��y"j�I�~�82��-�t����B�y
� �5"��]�?����ė3z�xE�"O*� P� $K�-acs��"O�P��l�=��A�;O�0\:"O�18�,Ѩ-�`Ӕ���\�(��"Of��g۔�����tΪ�"OV��$닢e5̙�O3T�!Y�"O��9��D�h��$�7�<-p�"O���4)��P��8G�8�XR"OB�����Θ�c�(_�2�4��"O�%�η<��7n��[����"OQ�7�M�K0F��ԊݎD��=;�"Oڨ0��`�`
Z"hfmr"OFy1�I�Bh�K�bϞOe��{f"O�;'d��>�&U�c�jB�Y"O I�#���h^�R��`���"ON���gN�TP$TS�J���	��"OlQ���+j�r�ɟe���""O,�xR
E&2�h�$z�� R"O$0�%c�U�R���< h�y!�"O~�a�G��l�,)��]1d`�%�T"O��'QsN��	ehS ](HW(�y�#'L���4Lߞ(��� ��y���a�������%~������y�L*���(���7�W(���y2"��Q�5Qeي�BQ�V���y�i/
�zY(%M�R�
���0�y�n�*�>��"Ɗ(R"Q	w�W2�y�,C��X�x�$��������yb/՞x�AyfoǄi��������y�F����sAB��2L�����y2���!�%�	"�D�fȕ�y��%��� FG�jp��G�y���M����!M;;1,�Y�E�y��O���kg&��/�nH���ybdQ�W����B5�$�S��ܩ�y"���z��R�������r,�yRN]'K�RV��:`���R�F��y"�Ge��;��&�z#c]�y��D�u� !b*�<$��ԫ��	��y�W�Or&pZ�K��B,�˔o�7�yr@��-d.9��+~i*��7 O��yR�:C��u�TގE�<�Ѕ(�y�$�3�)��lֲN��͐�`��y�%��|�p�EY�Ak� �&�y��il�A�8�����ܸ�y�"��)@�,z��@��Mۖ�)�yH�i@B9�P��?8g�ifdҟ�y2C�?+LR$c0��7��4.d�<	`
	
U�h���\�T��q���s�'���U��2f�*xP�$���N�B�	�Y"�|�&@�Y��sr��<"�jC�ɯR�aIb���<4ʀ
��hU
B�ɭCY 5$뎙u:
���FB�m��C�Ɋ(���Ӏ�M�[;�U���A�n��C�Ie֥`�kÚ=�8d��HBr��?����0{Id�K�2g�iZ�!SL��h���i*?�݆B�<`�O�Sάe�N^�<���95�F��f-7��Q#�X�<I0��=؄X91�M�<q ��P�Qi�<��!R�_�z�Q�I3/Su��|�<)'e�~@U���&~kA�[O�<q��E�fh"eq�'L����N�<q`	@�0���M�.wٞ�j��@Gx�%���A5��`��nĉr�a�*jh��^��� �ə�OɚE���۱�$iC"Ot��4��	V{��V��[�@}��"O�y�G�J���%�"���x�"O��YpB�D%r��'��4|�$�Ir"OXB�]�Y��ٙG�X��"O�M0!�.����G�:6G���"O��ؓ͌�J2�㱥��!�vࢧ"OjDӡm',���צC5��� q"O�l��ٮ)��]���P�1�b0�"ON0W�A&bT6���!�(!��"Ox����3]h���?s����"O|P����+e�h�Hba[*g`��vO�ԋU�D(c� �c��1$�1�64���#(r: �oY��V5A�e�cy2�	Q�'�!��Tt�-�U�L�ha��X	�'j�ՀaO� �<�bΘ�i[�'��u�b/�G��Ab냩�&�'�.�3X� CB�� J�)���'Y�qjM�4}r���P�~���	^�O����A������nˠ*�n��/O���3��|�O���Q +��IsM>z��!�c�'�1O��js�l4#��N��S""O�����Ț����b��{�x3�"OT���^	p:Ya#O�V�J�"O1��g1{�j���1T0�y�"O�TAᡖ�MZ~��Sm
?i�6��"OF�9�7g�6� 'j,/�>؉�"O~%�7� �_~��jbi�r�v<QP"O�py��D�^�R�9vH�(��4�r"O�t!U1M�1D
�#s��Q�"Oh傁�%�!�TFN�	��% "O�R����k�`b���!	���"Ozm�É�L�ՑBk�+^n��"O��=7m@�R3Ϙ3~} U
��'���i�HIu��p*"��:$Ƭ��:��K�O�OD^H���^3��KTC�/T��	�'vh��Q�*g�h\
�dF,%����'���N̪L�νR�!�6�P�'��u-�p���2"�(����'1�X�J�*h`݊�� b��#�'aak�̕�8K� �hD2u.Μ��'�6�"sD��'#����n�'��E���-�'Y��$��� �"H=�ܵ�� �&M��&�	w"M�u��&40ąȓ��4e��W-��Q��&q�th��h�� ���\�KK��A�!4�@E�ȓ Y�b�M�!�����)6� ���f~�& �5-��x ��9�*���`V'�yJ�%V<~TeAܔ8��m׆�y";f�( ��\0�~B5Ǌ��y�菏=+2�X&B����a)W1�y���4���D�������#���yr�C<����F�ф4��ܸ��[��y��S1,�P	��F)��P�����yr��{
���"��d��˫:'�'sў�>:����\Ԓ�l�4)���9F� D�zCHW�b�D���Ԉx���!D��s��^�(o(�7Mߪ#�tڤG:D��R���yRHʢ��;�\�Z�d9T�����eH��CH�6�:!"O�1�B�\��4�%f5a%,��d"OL�#�F�L����GOT�4rڴ��"Od��Bi�}�Zm""�N�(a�`��W��i�^!^ZY�"B`���/,D��  mI4b��Q��U*T(�=�"O�0JB	�n>� a�D������"O�I�� �F "�#�mX�CQR5b%"O�i���:�:Y�0��5ҝRB�Iv���a��'��T�У�46�"�m>D�\��M�j�4�S��R0�-�4�;D�`0&�]��K?C��L���"�!�d� �b�]!����тU�6!��n2�,��g� E�a����[�!�Č�4�$�93bQ�S���y�Y�!��څ+�H��Q$�3M�2(�� RN!�d�2���ɕ�Ě98쀙��j9!�d܈F�u�CN4|6��a�8w&ROPMB�D�[�j�1G���~I��"O�]��J�&�p@��*"1��ؠ"O�H3�+��R(�4�.+�~�B"OFIY���9q�c�-[����@d"O��j��U�h�d��&��R��A&"O� �d��e�~���@
�	�t	ҁ�I[�O=V����^��x�K����ig�գ�'s���eU:���C�_�\<EB�'d�8`���3j��m
�`)3�X�<!�(��d���zï�D~�9�G�K�<�� �1��e
�+�k�ћ��N�<�2b�[0f}�$
�p��s�N�O�'a�d�@��8�F얋nb�Xz�-�*2!�䇡]�] ��4UH�YY�+!4!���-�l�h�:	4�eK�;M!�
�{��UF�@�x+��_!�7>nP�G+LQѼ��� �^!� @��M���� ���^�!���;
� ��V�w�
Q����<�!�D�!����틏.j�����ت}%џHG�Ԇ�(d,R�.H1����JP�y��^�����͔Txt��CX��ybgL!Rc�զEL�=QrF��y�'ߩ,f�QS��7 ���֩	�yM�%S�m�.Ҭ�6�I�>�y/U�x"Fh��ƅU�)C$@[�y��M�	?�T���ݼ��Y�c� ���>�+O��#�+��� r0KC,H����Q #��H���E�f�s�(�p/W<KB�	{���CfʑP(J� +	hC�	5W�x��&S�N?�y��fF�+b�B�ɩ6�pkW+��u�X�@�,��B�	U+��c�/
>~�K��";{�C�	�:�i�4e �_�l	r�J��7|C��:~��iYt/��>�`�P�.�d��hO�"<ɧ �%>�h�CG�� a���!C��p�<�M2g�8��b�,s0�!��S�<I ޚ{	:b����Zt�B,�M�<�̈́���P��G�y�ҢD�<1T�=���r1�с)�f��d�u�<�PƂ	dVxA	Ќ����
�f_��8�'�ўp�<9��
\c)��-X����u�<�L
	ئ(�OL�����QI�L�<9w�	
qDh`Ŭ����F�^`�<Ye�)	�0B!fZ���Ր� �p�<q��(E4�!	�,S�ٺсRnx���'M�iK�O�8+��2#ʍ�M{r�z��7O��{bJC����哮y�
����'|����#�N��D���{�ҡ7D�\ aN�\���d��2���Y�@5D��!�C��*�M{��_,-�����4D�� �=9pm��V����e�֌s;\�J�"O�H���ќ|Жh���(s(�Pd"OX��Uf�m$���A�/)Hd�R"O�)d� 8-��h�2�TV
fE�"O��h6�3'Q�U`Ć^)�0"Ot�c"�,Q���1�,���"O�QHgc
+4"�zSJ>�v�	�"O�Y������;Ԯ
&���
3"O0�Ktd����퓷sc ��"O��B*sRr�;���rY��9��'�ў"~"ŌB0 � ��e$�Cr
�`�h�<��''ў�O�Rme�L�J��M:q��؀:
�'��O��vv�(� _(�4��'@�#vԀ>����PCV�~��	�'+�qѷDS:T�}���W@�a�'jݲB��Z3Tt�7��0zvTZ�'�!�¯�3)�j�:�)CI�J>����'|1�(@���]�-b���H��xV�8E{��I�>��`I̸%{�-��ዧA�bC䉟Ir���GW)v܁A��F�r*�B�	3<{:�2~��e+!�BI'�C䉃5�Z�s�i	���`� 1s�C�I%$�N(�E���|ʆ��S	A8�r����Od�lu�|2�铄v5�5$"�� �H���I\�?Јл(�{�Cg��-��@��5x�с�
��AI���W�� Ly.I��16�!�M�bg\�"��S�8
H}��6:�8�F�/��UJGFM2�X��LX���U����hc�F��|��ȓ�^@�d�J7sY��1%ێd��n���YÊ�3M�Ļc� }BhD��S�>� ��\s����	�[-fB�%�x�#�H��%��G�uX.B�I�&��0��F�"B����1~�.B�%%T�Y����0�n�(����(B�� e�l��U�N�DN��J��M0$B�	Fܜ�e�Q�z�KV,T�<�3"O@�4�Zz۸��aa�&Nʩ��'_!𤗚EzB�Z����.��i��̺	��)�'=��C,��s�EP�G�]�|�	�'�T�a�ubr�����+�����'�v]�a	 �&�̔�&�	7�6���'�������0@i�`��*�<��'K��㔂<'
���FT#K��A�'͚\��T��|1y��D�@0� C���c~���$0:�,� @�u�\�p��<�y���K�!2�.Os/�Abu�O��y"�O�r�X'��6V1&���'D�y�h�?�ZuR�A��}�x�a�Ũ�y�;y��Yx�-Wd�n(j�"���yr&�n�����L�[B����yraK��p�rM$[Ib%���?�?)���S�n�0q���#܊�:CL�gt�хȓk�ּ�v�Zk\���V�R��ȓ�d�t·�1b��Za@F'j���t�Ā	f+A�Q��`SeE�A��=��NsMid���6�"�\�DHͅȓ�,D��ˢx����eo�,�B�����<)�٨XX�l�b�X1�0P�TP��[��h�D2���s��W� ��1<O�"<ap@�&C#�$�f�Axx9B���D�<�b:uXl�16MV/m�sthI}�<  �4d����t���&��$�P�<��A�Z��iS5 �;DEQRk�b�<� ��c�
^bʬi��tFn]���'P1Oz�cwa��Q���R��$C2�
"Ol��eƚP�LJIЂ���'"O �	�� ������9Ɓ8v"O
����А |:"i�Z�hR"O���*�@Ҷ5�HG�Q�b�Su"O~|�!.]��Ig���6��X�p"O�E�UFJ�ca�x����ESشSD�'��ɹo�J�cG��m�}#��C,	D���?����~RV�ΣcQ�-1��])nD���<�s#.P}�Q(.H�^�J�'�s�<1���>��EK����|�����X�<�$�F�SR��N�q���EÆ^�<!Љ�8I�,H[G�W�m��	v��@�<yCiкB4(HGݹUM��C�c�<Q1��Jځ��.P!����bgUKy��'^l��!m����Cĝ<)�ԩX
�'�ȩ��K�J�x�kSg����0
�'��A�*�u�:HCs_���uJ	�'�h09��� g@|�s��6 $|(	�'�&hKT�ؽw�&=�ㄅD���'�Yr��;	V̘��A�n��'v���޺y�\dk�e�,+`�z��d)�*܉��BP�c�ڊb=�Q�ǜ|��)�?e��6l�?v�V�3���%0 �ȓDN\���T�_O�Y3�H�2$�R���N�6�RwC��t��&�@�-�Z4��V L�Y�ώ3tM���"d�"h�*)��"��M��FF�A�mF�tn���l��`�ՠ
��B2�Z��?i��0|��n��&�*�9b�P�n� ��/Ob�<�A�E�U	��ӷZ��bp��u�<��'���́$ ����: `PH�<ɠd��WE�IQ�.Zڈ�`��L�<ybBT�]�K�H��n��0� �o�<q��O?�	�r�h1da[d�\P�<�V�J6}����iX�=T��N�J��0=)���3:`��耨���[P�B�<��)؈%�p�lֻ~�l�GL�S�<	fGE$w����C��E�jX����Q�<I���)G�V؆�~�N9K�EN�<��+��s[f  �m�,�~���,Sp�<)A���JƤ�p��0�6P�3f�o�<���� !h̋k�
@� �'Jh�<���$����ǚ`��xy�_f���ϓp�꠸fNB�@.=�d���@��z�pD"��)p���c�%ʘ��ȓ*8�hCT���5����̛� ��	�ʓ� YX��ߗONLy��B'cRZB�I�H��b�cB~`J��dS~B�o�jQiƪ�K������Ϧ��0?9���X,�*$bZ3FX%��(ty���;�'!O�E1�E��8�ԍҏP;vՆȓY�Z0�A�F0�&I��/��cⲭ�ȓT� 3a녻N����H��
�4\��VJ٘�
S�91"�`��V~�@�ȓ���b�$q� =�ȓ��0z����P����u`;|��'Ma~����0KQ�I�mk�����yR��w�R=�!O�=bO�uQ�� �y¬w
�ĎG�r���ʘ��y�K	Ux 9S�K�\�i�@���ybE�E���pB	�-yǺ軳�W	�y��A�t�� A7�nt�M���ڪ�y
� �`A�K,2��!$M�l&,�"O��3C/��� �*�ԆOo*d0�"O�C�

�s�z��uI'S~��"O�Ks�4x�� ӑÏb)�Q"O�}��F�{HL�k�a	JP5X�"OD@���F4�Lq���_�9�"O�!�E�^�@+PAu)���6�yr��s�zE�U���h2,��y��,F5n���C��U����M���hOq������w=R�����6�p�S�"O���@�9`�P+bMS�o��J�"Oq#�����Ԍ�3���Su"O�<l[�[|j�0�ɿN�5�G"OLyjo�	x2�
C!��A "O�M{�
+Ez��`��5 ȼ"O���4�ςV����E��V���'���2w�Ё`>��uH�!>D�ACB�0D�p��)��U���a,5�{8p��'�,9"f����taf.կ*�>(��'m�X2��<e��僅�D�O�A��'.����e�nS�a�Q�U2Fϼ���'��=j��!�acB-+B�t���'��z���:�.�cQW�?t�
�'g�xj���V�J�k�̉�'���!�'�r]P� \�5��b��]��*AA�'W|�q��φ|���s�	�&�L�Q�<�ţ ���b1k��ЪCnAJ�<! �C(Q���J��͕I���O�<	���!+�u�"�E�
=�T�D/Hy��'zdJץ�(H&z��'�m�X���'#�����D�V�S��g������)��gəd��@��I��O
 H+"�1�yr��Q���F��L.���@�F,�yb'%�鳠B�C������ybK�.�Tx�F��h�4Y��@��yB́�wq����M��7���rS���'��D�D�ܥ��2s��"
<!�ϓ�O���t+ۢ{.�]C��c�u�T"OJ���%F� ��醃=`�	"O���d灝t d�s��n�EPA"O�`Y�Ȉ�&	�R'�RL�w"O=��*r6~�&K�5�:�Is"O�i�#�4Tw��H� ���)����;LO0}�s��8m����jId���rt��5�S��K-����Up��=*'�X�F��yR�Ɉ"���x��m<tH���P	nB�	�r�1�`Y���9�bܞg�^B�#}2���N!i��iq,I�xB�)c�8a1o�� �p��LE^B䉪r�J���?xϤ`��#5�C��;�2��b ��=�F(��J�)�C�;4��o����O�D��C�)6q�d�OY�b��[wA�;vHB��{�l��կѡcX\-��R%OxC��h���2��E�;�b%��DĽ�B�I�B�D�p`�^�(
am�E��B� C�̥,�6h�&J"/�-q�l(D��a1%WƜ��@�/%�2�o�Op�=E��YC��4S�I�#��� �
�I��3O�1� �ɇu��3 �X�`E����"O��p��#����fMM�ԹK�"OI��E(_��]�l�B�BUk�"O� �^Q�,��,%�<h��"OTMJ�o�R$�(@��}�ZUYa"O� t���W�ze��ˊ2"��)�"OF|�U�E�_Ĥ�bjڕa�� r�'z�	s�i>����8+���%�ҍ�&K_��yRiY|N�ӥ�|�,�a�a��y�+@A�@�i�#z�$�15����yR(շq^A�̊l���SK�6�y�	$��+�a*l������ן�?q
�'�� $n�[�*@����XL�y��'�d����Q- X0�ݭ �T�8�'��S�.�[�p�+Ů�{`��
�'�(��B��w$�Xel=q�L	��'g��z1	Q�{�*`��R�[7�Q�'N"Mx�$��5?"�+"3S[�9K�'ڴ1!5�,=� 4�0cA�Q+��I>�
�b)<	�$�[�v����M,%G�$��E{���ϕ3���'J�y� 
d�(�y��&/�� ��.����� ��C�I���RDB�E�����)�R�C�I���
��N�-��e�3�ҵh(�C�	�f~����&�UC7m�3efjC�I6�X扚�u:
��$ڀB��0`P5ҳ"ȌD|�s�+��OZB�Ƀ*�ٰ�Hڴ.���r���C�B䉎k?$0�w�� ���PƯ�8:��B��5X��Py�H
�%��D�K�&]��C�4�,!E�]�jGdh�2��(,�C�	o�t��l%5�N��"�� m�C�I'BѶ	�%(F�&�d��� ֚W[�C��*�(���晀=��G��+l��C��/�L8��#��T�H�8V����'�ڭ��0&d)���"UΈ��'��W��v���8�lݵz�b�:�'J����<�Ia�Y�'J4p��'BAӢ`� ��%�� �
���'���Ih�B�
�B��sRia�'�8��* XZHD���y� qϓ��$?�T �8�j�Y�@F�SAԵs2�}�<$Maٞ@��Ы{l�}�p��b�<Y�I�U�dm�E�+c~�ܚ �v�<�"���f� �:�<�*$g�o�<bK��S��8�f޸6,f�LS�<�gEE"��X���24a���_N�<YA�Ϸ`{�R7#í)pjqI��E�<Y�@�rE�W,X�D��Ck�<)��W�i��YzqŔ�aGh1�#D[�<���TO�~A@E�ֽdЭ���p�<9f�W&�����!����"/�r�<�d��(y��*L�V�4���n�<9�$�/L��p 0�7\=�g���?Ó/����R��33VIA6
ڧLd8��ȓ^z�UbL�1��B"S�ƅ�ȓR
�#1fJG��0�VG7/`.�ȓP6�E:p�H7E�,���
��po�ȓ6�$�"��MM(�F�7$�؆ȓ�N�!�<#�����$A4
�ȓ@����ƽ?�1��X���<'����c�b�(e'��l�tP�n�M"B�ɶ@������gy�T�a�RC�	>v����h����^��P�&"O���aNB�;��񱎗��tT��"O\�
�� �#�`�"˸s���P"OLL�UK�� E� �� <$��-�"O�Rģ��H>�p���2Z��3"O�e��#J�$\�ȵH�4�ʥb"O� ������"'q��'�4!g�y�S��D{���������ȏfx�T���ƺ�!�B"1Rњ�M;ZJ�a�"S!���i8��!��+F(��4oZ=�!��]#/sFp�B�$6A�y�iԎ!�!�UK�Xe��j�W��)�C��0C��'�a|��ˑu0#�eH)͜Mcc�	��y��G�dt����ʘ�$�!��&�'�y"�
P&��d��"X�sf���yb'@,�Ȍ83�C<Ji�kR��y�`�<y�xM�dF��~y8�E�/�y���G�4 ��� ��d�JV���y�C�$H}���A�0Z8xx-�)�yb��K�nhy��ү]�z5�T�"���hOq��I3�3��Hs��v��}�"O��Q�%[-⩁�JM">�8���"O�J�W�{mī�/��=���"Ot��V�l���SdBdߺ�ط"Or�K���4]��[u||�G"O��i�Oµf��UK�Й6^V���"O4�ᦈM�{�4�b�Q�h�4�'^�I<7V����ߗ�"dq!��j(�B�I�G�^�z�BVq��=D�>�B�IV=���n��1�Z�����Z�2C�	,D�!*Z�V9 A�;"��B�I�s���0,ҧII"��P�E>*�B��o�ִrf�]46�+ČO�
��B�I�P|���'��7	�i�.΢_BXB��x.��3��J0<����1�>��D{J?�B!4&7��6`�Ch�}�W+!D��K���Q��4�!d����?D���ea�D7����-�?�V�/>D������?��X:�!�=��:�=D��s��՟{0iF`�)������O��TG��'�x5�	H�vb��&$v:(���'�"���\�yQu)a�<��Ī�'g�$�V��]���㐁]�~Lĩ�':<q��.P(&�>�i3��o=�� �'����˰P��P�%�V�I�
�'��YCAՉ XՊ���T5hT�	�'�(]n-@����f��x�������<�y�d��(�9إgZW��Q`�V��y"��,`�R���d��?NX��#��y�c��@�[3K� �2�/G$�y��,'bF�`��Y'Q.hx Ej��y"�&;x�M��Oө��iT�Q*�y��)�
���M��,}��b�5�yR�"t���:"DD$��
��Z��y2��`pp�h#��
u�m������yBiU�4,�X��w𠣇�<��O�"~�0̏.~<��K�1C��۔�Y�<���VaǼ!�*\���� �X�<�w�B��(����yKt��Q��V�<9���5/���H�n���lوw>!��ª@��x@��j�"�����y%!��#`����w�%I���Q��<}!��E��5J�.��#tHK�k8\���v��� $m�h>��/�32��	�9D���!� L�z�	��&�1�tC�	�8�v�`��u3^�@�Y�+/�B䉌t(�AW��5aj�Y��e�B�ɷn�:%cĦ��)��IW��-Y_�B�	E��!>�H�Qؗ/\&B�	M��q�ȏ�7�r���M(DE�C�)� V�xw+&#kd (gj�� ���"O�M"��5I�[�H�n�XRD"O��`4a��;��@P1�5s�`"O������eZ�;GW<`�1"O�4�"�X��H�1�Jzi��!�[��F{��K���-���^�.���$ˌ@�!�D�n��}2��j��D�ݯ@�ўȇᓽ<(��s��*o��1r�G-�C�	3��
1&"l���@=�B�I9|���Ӌ
u$P�QoB�I�B�	 zĢ�-L�6{�T�ګ9�JC䉟7��%ڂj؋)Q����V@�B�	1LQ|�9�H�:/���iUARO���1�S�O���g#&��P�]r8���/�y���"!�`C�I"2f�U�J���yr�/~ ����Ƌ�WuR�t�Y-�yҊ�8XR��*�ONI�H�HD ���y�M1�)��;!�C� 1�yr��P� ��T',i�C$ɑ�ybL�)�"yP� Y��l
c	P*�y���A1Tqr�EwBDiBJ��y�c��&��2��F'Tݢ�a�!�y$��2���a�(�D�ŀ��&�y�K�1a6�*�:0�*j����y¡ڛ\؂y���n<5��9�ybd�#��1T]�	�1��P��y�+���ʹ�PO��}hv��J"��(�O�-�c
��LQ�D1�a�?5�QP�D,LO0aSGɴep���`��dN�d��"O��!>	yq�_��`�B$"O��{U�C�p!~|[��߈{�\���"O� ��gt�8f��Q"O> +G�]/�,K'�8i�J�"OD9�F���L����W"O�%R�(��"��������)��"O&�y���'�VyR�&I~^M c"O��q�d��	"�P�0vvp@�"Od�a�h.r����A�Pf:���"O��9����=DX�3��wc|�á"Oh#v�ɟ)�|i����f>^|{�"OL�*! �o̐�K��=�\$��"O�T���B6m���a`�do�8��'�ў"~�G!�;x=i��� .JT��j7�y� _w�Ig!шq�!�b�y�dZ�_�R��O x���b"���y����b��-�BJЁl�^1�b�^��yBǇ/�.��jw���ұ��"�yr��n$���[�s������yR"Ж&TaH� �l �T;��T�y�
`���r@��.a��%����%�yb$��F *C�����ׂ���y�B][ֈ(4%�jU�#mO�yRMI�'����ã�uZ�d�4ι�yrON)4D|��e��#�Q`D4�yBF�X���Q���J��#N �yB��UW�I���?	�T� �S�y�
O�3�̍��ˋ���R7.F��yR��#3�q��I�~��I�G2�y�of�YB��/Yg.)!��� `JB�ɂD���*uc�<k��� i��9�.B��&RV<��cAψL� u��Q�l�@C䉉���@n�,�J�
�#���=iÓ0�����J� d�!��sb"y��!P��m�+�R�"b�]�q��܄�S�? (�퉚_����g%Q3���a"O�i��k�7YbM$��0JG:�KD"OP�J�� �m�:}��̗:��m�"O��Xv �q��X�҄��7"OVt1@-����"+z���"O�ha`,�� U�`�6#Q?)�nP��"O|��D�Ľ4�ؘc�
�g�8��1"O���p+^ D���W��5{�F)"V"O^�Q-� {")�%%�jR�|r�"O�[�K*�t����������"OH�Z��9P��1jD�]�7�B�	�"O"I��e�'���J�b;��*a"O� �/�8�@	a�� 2Y�6"O�`�f(A�.^x�Dmڕ$/���T"O�!d`>4ܐѧLֆi�z�"O�d���R����7��yՂ�1b"O@|�̟�N}�H�Gۅ>*,-Z"OR�I� �1�^�昚z�^8�"O2��P��g`m)`F\Tz�$8�"O�R #�,�d]rVh�%WQ8�"O�0GHQzNn(!��N3�>��u"O��b�ԗ<T��hR0	$��qd"O�\���"*�i�eք�2�)�"ODaC���v��(�1
B.ݜh�t"Ol���``Jy"#hC/~�v��"O ���ʬ7���!%'�8�ЅB"O4�R�i��8�d (�5t��YY�*O��� ��6b��ԋՁYb�
�'�>�
�3H���B��8Fd�T�	�'�4*t���T0�����q�~Q�	�'����6��0q~��	�`Jm���p�'��-`�`P�EK2�ZS�L ozL:�'=b�8��.�$�z�I�rdh���'�����ݤ"��e-�o�|�
�'?��	@)܉���)u+�%W�ĬX�' �%1&� :p���"]�G�B=J
�')*�$��!���'��>��
�'6d��@�X�^�qV��3<�
�'�9�v��:�����h�%+���`�'�0,��h��*��/X���1�' ��E\�E�N�%C����)�'>���b
>|�晲R�>`?���'���u��#�H��q��#`S����'�^q1@W4�h���ij��'����ǠG������cd�u	�'��{Ѐӱ�RY`D`;`����'U�h(v�!+{R����HVjQ��'�A�WCG�e#N���`�>��t*	�'���1J��!$������@	�'x���Ɓųk 9� �)|� 0��'H9�%a�M�D�b��!�|�"O�J@�K�v��zD��(�B��"O�-�或�h\69���=qD\� b"Oj�Q�m��#��$�D�L6�Q�w"O�e1%�
x3�M�-H�p��J3"O�y��M�&�J��<N����"O��.�0@�
��_���ê�#9�!�<��0�w���%M��i!�N'K�!�$=W���2G�+u4,Qr�'Y�&�!�$]L�4<�$ީR��ۅҁ-�!�Ě#~DI���GM�Ii&a[6N�!�$UN�n����o1ΙȀ&��@�!�d�䵐T�Y1w^Y���
w`!�$�5"t�:s@��8>�=J���2R!�� �\��G,)�0���"�.<d��t"Ob��3#�:�>�p/��@���� "O����Yu_����X=[@�G"O��x�<5y2A2���@=����"OX���eӫE��0u/̄;���P�"O܅!��2@�����}�����"Oh��R%�W���*�b	,S���"E"Oh�CD$v.�C�a��Ҹ�""O#�H[v����p�'+�h0'"O����P�\����S;�Uh�"O*�C�~��PrQ��= v�� "ON����C�F���ťO�f̐�d"O�-‍�Y~�0ن�N���C "O2�)�-�<~x=;b�I�c�f9KA"O�t;��T�(�Z��sg�C��8A�"OX����y��}ʖL��x���"OT�x�e�+*h@�NN�D-�f"O�MP��ݵ;�b��ƅ(��U!�"O$\A��HF� "#&5�<��"O©Q����2�0���_��,�r"O$;bh�w �|��
�*y(�+�"O>�S�:w]4@�k�&p��a"O|\w��7S��#2�M�Kv kb"O��pq-h��%�Q ����"O|�UȊ0;��L��u���"O��K`e�qVb�w��=��Y�"Ol�{��\�u�(��$���u9�"O���R�N�T"*�%e��S���"O0 ��6.��k#E�H�B��"O��a�k�> h����+�P	�"O L�$(�SPR�a�)ީG�֬�"O�5��]"YQbǅ~Îe@"O@Sj6^�EC��D�t����w"O�sF�<֖`J��^�G ��"O��r1L�`q}r#g<
�H�9�"ODU嚈n��0�Α\�`j�"O8�c�پ! ��� :�ذ!�"O
%*�j��
��Р�P�Vܣ'"O:��B V�kS���`l�!`�4y�"O6ŰRh�$$���bCI!�E�"O����IߐmZ�cǱ.B�a"OHaQ��m��(�k_�$\Rb"O84���<s�������(�"O��;7���2��!�΍�lB"O�i3��ƪ�9x���$ �(A�"O��j��A6L����·w��уs"O�ЉSgG�j�4�vMR�,�ZB"O���HW�|�	�M�j��ə�"O&8�eՂ=���t���x *B"O"�/���2�fD�0���J�	!��ņD���Ő�ؐ�Ġ�:T!�;bn���gL��nMT����O!�!��˴t����͝-�h����}!�d��Nz.���јs!R��.H�0�!�$�6�t� �\�x��1d{!�$�e( D���f���c0Bɼxj!��E.=�P9���G}�����AN!�Şk�4*TΏ�]��Y�@�ݍ)L!�d�0�v�R�(*��8��mv��	�'���Quj��IU$M/����	�'�F����Շ�[$�0�&M�
�'>Ҙ9���)6��t��#HV����'x X��c�"J��hc�F7;_.�c�'4�̫���#�`0�b`��7{>m��� <<X"�S+�1�eGY�:4���"O��H��٦vl��c�ݐNڄ3�"O�!0�/����]ȅת�={�"ON	�ׅК	�;Q�́f���"O�񙇥P
x�h�%G*f�ހd"O&ā���0c8���hL�a���(�"OiQ�ɺ;�<pQm�:�NXHb"O�m(�h�%Z�fP-���Z�n.D�p�-�"e����
̋��}�d&D����L5M�x	��H�"���&D��Z`.��A:�P��b�R��0D�P�'D1xf~�kJ� �Fu��$D���Qi�
B۴�W
�=��0�E-D��j҈;\s65jEd�-P��`D�,D��K̦cE0�,N�7ό�5�*D�и�)��$�@��*�">@`��*D��HP��"s#��Uc��zl�� *D�t���L��$X��\\�t8FL'D��r���|�]A��π,Jx2A&D��AU  �Ds��
�N���f.D�A'��w��d*B��-��i�E�,D�������i��L�*��1�*D�@K&˅�Z^�a冞U�F�Zq�2D�\��@��Q ���	�p��./D�L��l��^���BF0�!�v�,D���C�W	~��(���!�e��*/D��r���W=�2@L�g�0 ���+D��r��?{Xx#��;ȋ��-D����"�hpCa'7����*D��ʣ&�&�9!��j�!ё�(D�8��.T2[M��z��*=��!�!4��x2�>(ɦ5"��)_bh�l@�<y�H��,5 ��"@L-�q��sx����@�^U���T'd�bjC�۞g�N���,�ΔQrE�,�pK�j��5,��?)���~�M��lP��rf*,���g��d�<�(�1<�H,�W��[��x��C�^8�dFzb�MC�m!��':h�<i��8�y�/�	�f�+r�K1ȓd��#�y"ӻWx4ѱѶu�Zt��í�0=)+O��$P�ԍ�h`d�u,) ��<���i�QZ8�F�	��x׫öDaqO�8FzJ~p��n�� (�i7��}�C�ZT�<A6̙�x��|r�k�h�S�L�W�'�ayr��
i��
uG�0%F�z�lO	�y�˔�(����@��.�t�0��y�oƚh�J�����,x!��5�y�W�&F��������熆��yb��z�T(P�}@�5��.��<1r�xR4O��a�j�H�/�V�x�K<D�$������a���z���s��8}��x�H�<���	ݕCQ�r�+�|��5��!���p�"�hEo��*�����A���-�S�O�p��Aq$ �醏�%���k�'m�vB
S5+���Pfr���JK��y2�� > ��aF�9N����CA��yr� +�,"A&�&;�t��[��y�͈�X�tȐ��$�X��,C���O�' 1�4��4�G1�F A��(X;~��`"O �`��ǳC�-Z�J�M1$I��'wў"~ڡ
�T�9�&k�2DFp���3�yRL�<�6XӠ�	K�`�����3�y�$�?���b���U�Z��ȒĨO�#6�X�'�Q��'>��*�aV`�<� �]��o_�w|�`�HևF��t	�"Op���M�,��i�%�cgN�'"O��ǧ՗KU���@�$�D11�"O�,��/�4"�B}"7��.z��M0f"O�:�H�$�8�0��v����g�'�Q���@
�(c���N�'6�jT�Ҧ%D�h��J�.q�>�I<:�%�%�d=�S�y�XT��e�~4��D�
,H�ȓ�z��C�L*J�ԡ{ a?_���ȓY<���J
Ӏ	�QǙ=;�m��]�:z4CI�%hX�cB矢�������M�o� W�J�ق&�p��(0wa��y�BR�>�@�!IHgQ�=I&���y�%Q�Q�����Ϫ`.��ڵ/R5���8�S�OlB�rTA�F9&��C8@�L��'ݠ��rD�<
/>�r�@޹4F,�1�'ڈ9[1�ȭ�9�f&,�z��'4�b�6f�AƇ�B'��P+UE�<!b	 ,�0�FM�#S�N-I��PK�<	գC-h�u��2���+�ǗIH<�R�8ֲ@�A�ѡv�|�G��'�T��	�!�r��'Y�%�Ĩ'	��M$B䉤Sd�1(���<ل}�"�@.@B�IYIl��6�M,BL�i�-��*����$�y< ��g��.k�4!B∔<Z�a��	y?���,������C5�����6 � ���k��tW�'3�~Ȋ3c�89�ل�?,&��Ň�
?��*0B�W�������?E��O��[�D��ԝ�֨��B�̙�"O�<�2��r�p[�}�Hxc"Ox��f"͋���@�Ci�h<�"O8T�� � ',��G`vX�h`�34��	��F�t�ih4�C=;��蠵�6LO��|1�-J-eFꀰ�-�g���pJ3D���D�	�>��q�4������+���OO��S�3�M�m�B��bΖD鄉8���81!��V+J�`��GCӚ�̜1@D�1i,�=E��'Ctk��/�}�C��
�4���'H#��	8Iu`���f�kHT�'�9@�lԵ���y�gМ|��c�'�j0R�
X>r�X���?Ik�4z�'��T0�h�4q���P�@ϢA�'Yў�}R�@ģ0=�@�Յ�$���a2��@�<��MP.uX���q��SrP����C�<��D�;K2(`��@�qr؃DQ�<�Mp�Ԉ�� O-Zٓ".�A�<��ſȂA� �K��Ћ�E�}�d6�O� 9!m��(���ItEeK�KQp���+�8OȽye ����k'�ւ�F�#�"Ofh���c�"i���F�|F25���Io�Odܡh0LC�q�D@fgG��58�'�\�)i� >D�C ˴�r2�'�K%��Ut���n�|���'�1��O�/�B([��'yN��ɍ}b�)�I�"%�L�`�/S!<��S�P�;�!�$\-P�&hj��H��t�2�MW��1Or���E�^�ĭیx��Uꄍ�k�!�d{��آ� ]�6��Zs�#]T4��m D����]�ji��qĚ�2X�<�*>}b��h�'>:��w�tV��G̉j�R�r�C?$�4ٱ� }I��6��i�Azǉ/?���NRya���?#���Z�B��v����΅�g2�x���M��C䉢ctZ�s���iyѧ��"M�C�)� �1�e��$_��:�N8g��M�Q"O�$����4�νH��{���:��',��b���v0����0o@PCtȆ��y��'��F�_	o��$c�a�8���D��O�D��ۢG��K��
T ���"O���O��%����ZĠÕ"O��x�D�R�^����Y':`�#"O� �B�dxt���E�rw�� "O��qI�	Kt5Ii@(k�1��"Ot��_��fW7�Ā���u�<�u���]1@��UK1ynjx���w�<a�M��_�$(�Ͱ]w8 w�Ru�<��ܨQ�XCF�T�%O��kc#t���hO�'0��p�l��8g�5RcjDk�ZP��:�*�أ	�Z��9�Ƿ;��$�>1 n)<O��`#� �Ab��&k��e	bQ����H�*�P�A�+�|�#�t�Tg"O��SM�?5��'AX�z7j��0����	.O�p�5F϶ 4���``�9>&��d%�	
p��i� �{=^��0��!�PC�<�H��'��8j>[ф�0yF,C�	�t�L`Р�Ǡ*}�  �?�C�I� &"E��+T��A%);zC䉯�R!J\
�`r׀��@���"O
�ѡ!�7	*�e�
��6�KB�i�ў"~n��g[Rm�b�I:w�đ�j��)��B�	 ����� 7hrFض�A�5��꓃p?I�
Q�L�Q��(�daQ4��X�<A�+?F��pH��>���4lR@�<����Xڼu
D!΁S��`���[�<��O��'�"~@̱N2DT%#�D����w�<y�aB�]�l������a�p�_�'K�y�� �R幡.R��B(����y��1h�7)�'����i���E��>�H����R�"m"�-�%Q׶M�ȓg$D@q��G~�&�Ĩ6d������W�RX�WL(|c(�����)�5JL�}�tuz�+'f�:݅ȓ^�\����-H��)���84����ȓǤ�y1*�_�N�a�I�%���.��Uɖ��=-(�1�ǡ0ϼ�ȓiȊ�eI.a*�x�F��V8,I��cRuS����,�m����7��)�ȓ ��2Rf�,h[�,��K�ņȓ
f��1f�V.��h�\X�ȓ�Eځ�ƙ�䐛B�ča��,�ȓA��Py�b�b�^٨�䞕Gt�y�ȓO�z]��&��Sǲk��˨T��=?�-i��#Z��Z�G���4�ȓd_н�p�ܑu�X��E�C=_� �ȓ=�V����Om��xbQ�ҷ�؅�rd=�I�+pd�����(�ȓ��l��BB�e���`�ˋS&��ȓ5G֘����q)"�F+�~�V�� <Hi�.��oA�"��\>EO�͆ȓ�Nٸ��0`LxM�FA���"�ȓ'h�<(4+U2S)����$�ȓ5A蜳P��?��8` �V�@e��u�x��f�,b�!X���.xPx��)��l+%h�딋'RɆȓ,;���ϙ�FH2�K�����D��ƚ�b��_�k����6�פiEd ��ul���Z�.B�Ѡ�"^~���ȓ&r�P�*I�~&n`�g��F����S�? ���5�1R"V�c�.ѹ"O�[I�:\���� K�
4�xH
"Ob�"Q�XNE�9�,זb)��a�"O X�r��R������<vT����C�+��P��'	�3�dY�E%���l\���8�'E(�)�	2�i藯 Q��'��I�4,QDj��P5&�=h��@��'�"�Y���<�P�A$��/jz81j�'�:	
��ٝPr�d���G�o�.��	�'bh4i@��L�lQZ/��e]���'Ǭ����Y�FIN�j%L� �L�9�'N1 ��>W����4��=��s�'u�S�I`W^���w�n ��'�`hR�I������#l���P�'4"̓d)ڏrޚ��CG�=`vN��
�'��d��*S8N�����b�^u8�'�
��(��*|�!E+ǚXa:T(�'�N���܆>�$`���&�R� �'v��	%C�_�*]�3+�)�X���'��l��Fc��)3	� �a)�'?(��A� ��0Qs)��NҮ!#�'�Z����6K���`D7F��H��'��H��D�
�$��7*[�vWH�I�'3]�F(�)M�x�G�,�ڀ0	�' �`�iK�|�>8��]ag��P	�'�"����W�?�|�
&M�1g�.�[�'��|j�����(Q�%��V%b(�
�'�H�2!�օ=�r�G%Ar����'�Фl�>!�R�i�V6?�@mR�'7BeHs`�|.�8Ph�&Z,��	�'Ut��E!��P��aA7Q��'AX���^�m^�A@��P�:��'{���f́ 󾈰�떩V+�!��'��H�� ��!H�h���-�vP�'$�q�s
�>V8t��S��t*	�'�ބ��
����#�X}�L��'�b-ʓl�<I���RW:i	.i(
�'&Tj�*������AU�P		�' \
��*.����J`t��'Z��H�4:��%!�dBR\ ��'+B�62�TҤ+J�K�>)�'������+b(;���$E�0�'�tɚ�c�7CU �� 2����'vbp����T�y�
B-ŦE��'�:�/�2t����c .W����'V�`$�_�x��(�2K�8���:�'2E&��"�,HB�'��]�qP�'��i��"�6{Rε�Ď� d p�'֦5��&T�6[|(���<&�0�'>&�����( �<]��O����'_��!T��,���r�ȷR�3�'�4![�f�>�R(1��̰A�:���'����TD,-�@�!�+T,�<�'��+ �~��1f�ÇU�����' >�	u�/Y�D�1�KN�H�4�i�'0J5]��+t���El�x+�'#ʙR�kV�,`��8�"�'?H���	�'���G.F�(�RC*(,B��:�'E88����-B��1�M��䶱��'->����yGLjBIB�z���'JT������j,SP*
�\*`�'��D��bR/.�����/����
�'�L��K�B5��(��/�>�`
�'�0�VfÕC�:�a�;k���Z�+��q ��'�� T��ƎM��5#fIԖE���d"ON���Fٛp�e�i�r�)���0�$��(PCD�>E�T�¼�#C�S}.���ŝ��y
��X:B��炄uC�}�r�O�I��p���O�b���z�\&>c�,�r��5V�(�/1R�r(�Rj.�O�������RupjL+$@9E�L�L"��`s���}ؔb"�O�5���U	�س�Y�8����I+PwB�j�`K�h�Q��Ai��M�L�����V�!�(a�����yr�
1lB�����sZ�Pv �$�y�f�P�yg��a �]�E�
0n@#}Jw%իYT��C�
^�V� b6Ui�<�,X8^�֝Qt�O2l�N\�]�<;F�4wb����ۥ^|�җ�?!�����k7|��ǐn�vL��d�58�}�$�:����C�	��K�ӹ6#<��b� )��U� �8'h4�SC�(_)az�
�*p`��1c.X�څ"��W4�hO��bQo
��n�xEk�>r�ĕ��M)��� ��W�S���9��ЍXۼ��dd4D�H���q+<e���Z��E@s@�OX�1�"S�zF�����1
a�7.��r.8�?�*�$�$�>u�%�0v����A�J�<��E��oy�8y1
�N҄J�*��iTDU�V'���4[ADL�c�OOX�j�� J,LH���M3+���
Q���}B���)�B�p^(,85χ��,�+ �׈v�N�i'�C�W�hH*�9 �azB-O�jj$n	�Y��t����8�(Oh��p�U,L�x)2��\��T�6�G:,\���
b!T���g�jԌ��bD�y2o��-��!��V2yJf�_� ����	Qq)nP �P�a�i9R�Q;.��)����b��d��!�j]����/�vA�ȓ�J��C֐��$S�G'� �� h=?n١O36�l	�NC\�Yw?p�a�y
ʴ9�ԝ�����Z���ic�P=�0?�rȞ�RW�����PlT`��L�C�UY�+;�1�F��e�� ���<�Hx3x��gI��+��p����T�'�"�W��*{����BL�i!�Tѷ��@&),1`�oL7@��2��14��5��58��f�(���j��Ĺ�H�5�H���U�̹ʠg�ܺ3���ZS�&XP��A w�蒖���y2��[�Ypucـ<�f\�6	R/:<V9�5@�T2���R5:e���^�s�H�$�0
2��(6�2$8�hKJ+by��-�O�lk��H�eʾ��e�I��f)!�Lgq���blʚ[:��;���1%�6nAO<��}BO�2{g�P��\�)���%.���O�<����K�5��A�;Z�8�oݭ�\�7�j���C�@A̇�N���'�a{�#�2#M�X"�G�XZS��U�~ҭ 0�ܐ�X+�v���ِ'��Ig>��'�ug���H$S1ǃ1ڞ�AW��yB����!j��Y�
]X��BC]8#��B���wɚq�pį/>ڑR/���Y�x�Ӽ��g�,	�Di����;�	�ŉ�i��x
J��O���K�E��VC��W ȴlK��+��
:6]�pDZ?p�'�y��5ʓvd�h�qhX�� ��o%	�4�E}bF'���j1� A̧e1:����J4�L�sf�&a*����~b�'�� �baޞ/p0�"+3G9(�S�'���H�cYZ̜=�O�ӕ����O�h�4�S�N������k��Y�"O��+�M1##LE;���)�Z�ag�xb�M�(V��B��z��㞤�Ӻ;��q�t���֭o�1��g�s��8+!�4'�p���蛭 �B$�,��j�-)i����<a���yb�!rz|X�-A�zy�$���yR��+*ԫ�e�V$QZA��y��O2���Z���'�4O����2\����>ٛ'�Z�1KȸOf�m�Ï�73|u��'�z��T�N�m���#��"���s�'�����S�o�|����;f�lM�b��[��B�2@(5�Q�pRXAsL�p��	3$�~��(U�  8�lP'X�u�����p>I��#?�t��7�����fi�Q�$��W�<���Ϣ2$L��u��r14�#N�Y�<Q7���&x�[SF��Gh���o�P�<�5[�^�8��Y�wntѐ,�e�<ɡ!=���!b�/Z� e,�g�<I�� =&!v%U#�|8y}")px�(A7i��z�
� f!ږ;\ʝ��:D�l��)�2m����
���2.-D�� T��E�[{�V��#��D�����"O����V�m����1�0f� ;C"O؊"%Vm� ���60��k1�Ol������d!Sk&�F��c�C�	?|e��l"�ΰ�G�B�W��eb��$�9&~��w-	x_�0/F2u�џ�E��h��mu��v�<�8a2֤�Z����s�9��#	/�x�H�:l��'��LpI>��4pn�bs%�E��� �ǉ6a��X�ȓ�40�%�,~�d5ز��-p�5�'���� K�r��.��!�S�]PF���%�Q��R'�0v���=A�%��P�`e� �2�O�q�1�O2x�V��2]� �1\�d���[��~}*��&n�G��nAQSH��X�N�Z�g��=�Ql�-)n ��R��(WN����O����JA�=XW����3`>@��V4a��Ѡ�'� h�΄�'��z�,U�mhX��ռy��RD�ґ����I�R��͘5�*F3&q�٪���z�+X�]���	��k��6R�^��Q��}���s���@�@��I�0eRňU����"f�\CU��*�뒀	sp�q�[.f��E$�K�T�69�@��ny2�0�'(z��T�?3z�LK�*C��Ey�-b��$�<?n�3���FC!�&ȡ�m��+{�y��Ɲ,l0ʓ Ơ�9���}��O���qT�����@��e;�\�F���Nݺ��J+(��;㉴�?E�$M\/���!��a��	` I>D#����4,Ƥ1V����	�Pi�PL�9iC��IgaH��l%�0�����$�w�t�!.�Qm�pS���9jG��a/OB�aRLعr�����C�G
�"D���p>9DK�wiP5#��]�8ǚDR��|����f��b��,��lI� �:���i��".O�"}1�E)K�@1�������%�C�'X)(A`�(H�L-�sb� ��O�����>dF�Q�)�2�|<*��>�`�`�Xt���}��Ǻ���l�rs҄A�;kLz��� �,Œ=g�MEA���ړ��i�6戬]�Xڃ朹s��es��6ha�B��>T,�P�%�;�L-��J�A����R�Z���hT2:��\
����8���	�"Bx{�GƇ-�I�w���b��$��x��������M��cX�1��ݙ`��z��y�u�R1o>Q�G��'$���Ӯr�Ց"�������a�WRP`���Q�O�BHTJCe1�����F�m����'�6 ��ɝ� �C���F�%y��'�ȱ�C8rc��yL�0E��'�zY��B@�\A�I���K)i�ܠ*�'j A�#)�2�܄¢�M�v��9y�=�\PA�I̪/�����=��8S�ۮGYЍ��"zJ�{��]�>&�H�ǄDԦ�1��5v�VT�r�Z�m �m����c�$��S��?I����*�z � -�De��W}�,�8��� �X;#}��f��D�uL[$Jcj�S�s~B��v~��'��9kw��f�`$�$�K%8��@�)�2t�� x&�|��9O��3�����uA%H�I*�Q3"O
�م����u t(�,��S�O�Ƞ�!�0>!whW�RD �`��Qq�iBs΄C�<	P�?Lթ�GL�C�ҁ�p�<)"�Q(v��G�u8d�Ʉ$�h�<�ȕ%p�Cv�Ş!a&�׊M�<	w`�{@jD�D��X��vHE�<�掍�,���a�T�i,U[��
[�<�)�?!�L���־�.\{���S�<qGZ��P�!���=��1��\E�<�Vo��E�p��#^�Ɯ-!�B��Yi����ՙD�Qy��#l��C�I�`��Ѣm�}ڡ�SO�${�C䉄��� Ћ�'.r����gJ�n�hC�ɞ_&\����\ VA@��Q5�C�ɦ�8�
��Z,UTH���'�&$W�B��q/���֯��,�x���L���B�$�0�@qU��I���	OV�B�dZ0QBf�gq��˓��01BB�I2Fe.�q�H�*�ԕ1�E˝-�B䉩[���Ĥ�)i��%�T	�)q�C�	�*�d8�Ɩ,&F�)�fĈy��B�Id|F�� I��������� >TB�)� hYYE�Ε@�L}+A�I2	�Pp�T"O��`�ND+.DZݑ��*=��tz�"O���։�k�R��QlA%7�����"Od���ِL��+����@��y�"O�<��(58-�B0R�t���"O��!3H�D(�	7A�1E�p�ѐ"OT���瓓-(ZH)5��t8q�r"O.}��oIJ��d��_�H�"O��	�*�V����n�
]��J#"O�,㱈ڞs�hv�&y	�S"O.��'D��)��k��Ǆm�U"O�*2���x��p	�*U�Xޔ"�"O�I±i����ye	�Dj�"Od��֥��~C`Q��fQ�^���"O<���n�	v~(+��¨]�4*�"O	�&�X�(�.1�ȃ�O���i�"Ot��L(#JH�a���{w) V"O��H�DA(zo�Lx�#+uzl�qQ"O�P���*%��AZ� |����"O���B��X3�$��5e���5"OR������)�Qj�k6�
�"O��S&�>�I���v����"O�ف�A��_�4��c�3R�\��$"O<����Q������Ȧ4����"O�9�$	_$l�V.@�9rHt"O:!@��<:��YS�I#tj��r"O:@�����__�q���XN�h#"O ���\�=LV\�5�ŗg9f�X�"O���G+�]V�d�2�D%�u "OX�,��;ʾ�� ��29(���"O
�tK�2�H�Do��Z���Ä"O��*��9,3�1��H�y�A3"OBl�EcŀL:ʀ���F�8���"O  Imαr��s�cJ�m�<d�P"O��qB�_�z�\ɡP��-}6��9p"O((��LQ	-�Ѓn�[����V"O�9P��1p��P����A-T�Y5"O��@��<m�`u��$ktaE"O4�y1LXc(�J�"D���2�"O 0��&BA��H���ɗ���XA"OYjf��Txh�q�ם<����"O��Ȉ/6:�MCT͟�P9�=��"O"��5��.�:��!�7��ђ"O�Z eN�<M��
�`�A"O��j��8�A��؆�]�g"Or��w�0`D�x�I�	瀴��"OV�"��I-d�Ea�ǃ��p"OR�a����I��I�g�.��"O�}����(NE`�'�7.� u��"O����� |����F�.wȍ�d"O��e�N�uɞh�DI6Z����1"O�@SM&ب�
Ad��5�>� �"O~��%V����c��i�T�H"O��X(M���ktH܆3Ŏ�x�"Ob���0zPi�D'Y�ZT��b"O%��B�9>�Qc��C'����"O�xI�*Q_��|�g���~Jܙ�"Oz}�1F��6��PwI�N�ޠ�""O~�H��8%�b�ǂ/B�RU�b"O0�Ra��%5,��D	�$]l"Or�yV/�-�D��F�I��ԣ�"O�4
թ�#�:z��nh���"Or��%��o"�Ĉ��t�zY�#"OB�x�OX
]�x\a�I�4~�2��"O� �Y9g��9<�P�t��+E�xѰ�"O&@pe��=� "�.ޯd�z�cU"O��Q���tw�I��,G�0� F"O���	��Pƺ	A#*��6�B���"O؈��La!��0�ս#���1""OApbQ�I��,��^�
��V"O��%ϕ#�lPH�H�c��-�"O��s�iY4=$�x� ř��١"O�tZ�+���:� �e�#RB��"O\Y'�O�P���#UA:x��4��"Ov���&4�"�Z�(c\�	�"O&���c�+x���2� AH�^���"O�k� ʗ�J|� �յ�����ɛy��,��铐Ifl@[�f�#:u�&�&qM@B��%f(����=}����*fv6�C�`�!Ӗ�/��s�؝Pu�t����3&[�1jZ�X2"O>�i�-.h_ZcP�B3WjY���OrIӲ��!��Zӓ2��QC�GT8
v���'S�F<�y��N'
� G��t�\�+���D�T�6��5H�p�"O��W���?;xˆ��A�!�V�>��M�9�
�SBM� r���''§%W~9D"PP��6��:�h��F#	��L\n�d(�$g�Y�.Tk�Q�:��U�6�Lp^��eo�u�g̓4����Żz7��fȆRY���	�5��q�Ĉ�v(2	C��� �[��dI��y��S!4h(�Y���y����B�X�p���V������&�`Ol1�!�µ1`\�Swkߑ �@ � ��/7w)�6OU�y",JozM�5�ǟ$������P8���u�4��nZ�B�V���D\Qv#|"W���_�.� ��O�r�e��K�<��
\6h�8Y�1��x�\$ e�\�y��q��,�A�I���D�U*�Y$?�pqe�oP�&�D'z��aq�>�O�e:��V�B��Yi��Är�:\SA�G�UK�Z56P�C���=��$�#�1��� 9v%@ר\�'���f��=��	4@ܡ^v$1��C���Vd��1LA�#n���4��q���i �vfޭ�U,��Q̖��'�Ѕ)w�W��^R�]�0s�D��G����֚5Dr �F���y�@��q�2c�<&�ܬ���%4l�����0�*�s�+MY2�x"K|�>9�`�3�ެhw�ľ�Rs�Z���0�&H�HK���&N 1��	����e�m���l� 3 @Θ�P���)Js�����,fɬ-ZQ�]�d���>�tG�|f��2�[���a����\w!"5a�'W�*�Ӄ㚞m �!�'M�8sd�;:r>�Q�ޚԾ9�'q���3��-�ڈ��M%[��)"�S3��DX!勄f?`$X+�����'�y
1o�M����lҒ ��C��&�ܜ!�Č.�>i�L�/��3��8i�D:#�X7

�b�*��4����d�1=������=+�(�@� ��ҵ���)3Rɣ��
u��I�v[��H"腇6�0����d�D}�O� �JP(Ï�y̧'�Z���%7��x�杘�0�ȓ~�X�p�`Y��.4���G9b�a�� -AY6$<�ҧh�.��g+V��m�'�U>LC�e�T"O8���e�60�z��.j�Hu�xRM	�_;�,�0�'F����\� �V쓀lMz�����
}Bɉ��`��B�4~ �1�ͱI.C�	!IYL| %�Ϲ9����ۙI,6C�	YI�l�"L^<� �KB��'V�B�ɇM=����}��c����
�'^����l*�$Z�O
cQ�X	�'���#盯�����̖n��5h	�'	�W�I�,Y,r��U�a�,��'ؠ�B�R�$���(sF�<^'T4!�'7�K�*��T܀<�r�^�V��
�'b�]gK��f!�mr�R!T��9��'] IڧÕ-��	`��=w8�)�'��ћ#'�f���r�aԦE�t�
�'�F�x�F�*�F�2F��2a�@J
��� <���LS��t)���؂n<��2t"O�Ų�(Ԧc�
9��@�my["O���d��{L�Q�#$�,s�����"O�y{��U) �z���D�X:"O.	�R�aڶ�4L�`���"O��EB�Y��B�Yk�$J"O���H� RA��7ay���"O��!�mĪ|��4��dL�a�)��"O�ݡ!��~���2�-�=�$"O\����" �>���OSt�P�
�"O��dퟩXL`aT��Z�
	{�"O@-�$�$g�2`{��W"@Ȗ���'��H	c� ���(��-jU����'��E�G!ϵ"�
����12Z<��.O�L:����ʒOQ>qhu�L9$�D�7+Y�if���/ړ>^�)s��	 ���B��Į\�~�J�`�U8�LZa`�A���x���b�;!����'��@�#D�'O��5A$�R9�8�zܴH}��ڴ�հ$��M�g���?ub��_�Kx|P�`iςg��t��6Z��)�'���(����>_b G� �fk�h�bE�fh���'�LР�NU�t"��o��j��U�Ȉ�tU��.�1KW�ǆ%�6e�I�q��|B�4#���CK1����OG�`����d�αR�� 㴣Ɋi�~�[�ڝI� �[��G�# /R�k"���2��M
D��$�(O�Xʥ� %\��@1����L��eϼf�q��M�)���c�#HTy�G2}� "�όN���Ū9���E-�4K�T�1 G�Q/X���*܌V��Uq�L�xL�)§I�P�8���b\�(�'��V��� �����If%ɓ��?	0�\�����	(�x���`�8����:,ȡ���V�."�kܖ���c��/���ﶍֆ��obi(F �=�t��g�'�`8����i喝��h�L
��3�5^r>I[4C��_���ᔀ
8�`E�U'ӵD2�	B�O�6e��5x]��*I�HѢ��䐭x�8y�tF��{Z�)�
)�� t���hpHC�N@�F��;i��'���g,R�u֬��OVq�al�&v��JZ�JnsqL���|L�0⇏s�����O�>K�1[�VP�2��K���2�V,Zv̢e-Ee<ATE�i��;i@obh��� ����8 �
�1�f�N���	4f&4�[3@�O�ԨG�]�+�����s,�0b	5�M+��42��a��-3�QH�<�`�]
#�n��lOG>53��_��g���SAW9C�#}:7�̈́+��ӡ��%�"t"�OJW�<y���u�����j�N5���9E�4i �'�z:��h��d�7�ఊAJ�h|�0��FH6L�!�d�&�@���J��d�d��Fx2�Ċ�p�K�F؞�+��ٗkf�s�#8N�bȓ��8|O��Ti>lw��;ݴL�T�{��C2�hr@�+� ��oB"x��,@��p`j�#����?�@dyي\�L!�'K��m�t�plu�6�$�؇��)h'N��Q��4����/Z��;1N�t�́M>E��'���d�U� �FāDMS74_�A��'TU�����Ȥ�'���!�J�'iX�0gf��t:C��B-��R�̡ U	�@ȄB�IC����T(�����H�Q��B�I�(n��C�ӛ����J�?Y�0C䉡y��4S��OxG�uz���g�C�ɔ#��I{D@o��i��ݡX�~C�I�$L���V�/��ѷ�gvB��+s�ؙ�w�F�Nв�c�+YB�=A\J���	V&q�I[` �9m�B䉢!l�iEm��7P�mk��Jn�B�ɡ�\A��'O,h��hS+.C�	�,�r�A7�[s^���V��"��C��C�HAP@nI�i���%�<7_�C�I/i�~@!F&�2H�������7jC䉩{��e�ҬA�P�f(ҥa%8&<C��,��n�����(F�Z��B�	�zC�cS�0<�V\ �˘�4��B�	�
Ts�̖(;� ��d�B�)� ���(#9�Ƭa�iڜ��`�"O(L{# �zp�ЏC�I��)ڷ"O&��jޘ	�<=�뀄4�P�*�"Ob�kw�z�: P�Tj���"Ot�����F�h���͂k�l��"OF)��їc�A�lLgH���%"O8���+@�V儴���$��"O�ؙ��1I2� ����]�Ƶ�"O��L7�8��&�zp�"Ob$)S���	����P��D��"O���� �$�6u��H`��Ȅ"O��P�([�̅�sf�K��\�s��b��ʵ�'	E��c#h��ШŊEo����	�'�f�с �+�P9���n����'`� G$�Ff@e�*zTp��'؜B�������r7�ԋ`�@�0�'5a�#��r�������]�j8�'�,i���b�iY�ʆ$%  ��y��Ƥ�O1�Ve� ���fyj7��!<V$8��OJ'�;�1O�>xer\w
éɲ�� Pg����@���S�O�*�s [�4����ԉ,���H���0:��O��@��ɵ|bC���+ZV�u�O8y��� ��M�`U��#��G~>���V���	��'e�L���}gP��� �
"J��pB6One�g&>�(��O~z�jD��)Qh�˲�.�J|z�'�>��Z�h����)���𩋨�.!���'BW�}Rb�_��C��$0��T�
;OK��S�O�$��-�"Lb2���l�<P�mҩ\���""!����)�'�u7���O���d��1jW��,!H��J�>�䓡0|Z�o�9 ,931 �_�6��JU����'Z���	�@T`�����_���C�ާ"����,�F���j�<���d�J�8
çk�݈c���.�P���Eȃz� ����~p���V&.Cҧh��5��3����iP��*�ᜡQ"\d�'�ʚZ��S�OU�eHƪD�yn0����*����G�d�H��O�����OZ)�E[�'��(��`ћ�t���Ղ��7�����O)�e:�e�����b�	 ۾�:�'jTȘ�C������B'����y��'���yu�AJ��(��-��'}nѱs(Q�9?���+}�q��'
��0��7E֦�i��>	%���	�'J�&m�0G;:t�D
>����'`>0�c���$ry�U䋃�b`��'}�!ʇ��"���9f�ѿk(X��'���'��#����`��\pA�'��j���4H��uj�a�: ��L��'t��j]}P܀�/|o�ܒ�'�y��(<I4a��CݷG\��'`0�(3��X�
�3J袤�
�'����vLN0N�ׂ��C���J�'��Ԣ�O�`�'�-.��|��'���e�O/#f�Iٶ�ߚ:�
�
�'�D�i�F�v8-vhY����+�'���Ti��o��шʐ���'�H �����&���ûN���	�'�B�#��?\|�س�6X;�J�'
xĺ�Ñ�r]���h�%�ab�'ˌ�v��+�$ �cf�
F��J�'#P���U�����	d�����'�T��%B�\|�I�f��\!	�'�@pru�ˋ^&�)H�� �N�HH��'*Z-����0B_��IS)�;L�F"Of��E�?���I�E���8t"O�,;1 ��{�ܹBP��urpвG"O�0@�&k������Z�� �"O��@ 	¶�\Q푉X�,3%"O� �ŅĢR���,�=XH�`�"O� n��׃�_,tY�LF�IE��	�"O(y9 �ۋ0]X��Db01T��B�"O�9�L�Z���2��w:���"Onu@"�׳8��N�j7�-��"O^�
��~���/O+Ҩ�Iq"O���O�4rpD�k��M#]���)�"O�E*�o;F�%Q���X��"O E���
 %�PRNZ$r<��"O�t��K3@�сҍ�R�.8�"O!s��<�6A	�*�X�|3r"O�� ���ڲ�*�Y>2�0`"O�aqH�k>5�F�M�N�"ON�ٱ,�h�Zs�Y�<�2I[�"OubrFP=c ���fM܊ޞ�#"O\�QP�ݳI ���KB��6H"Oh1���#�(����;�]�"OX����/p��
ӉCX�0��"O(��S�-M��
�
�\���"O7�Ֆ<>���kΙSa�M��$D�k6��9�6��t-�=@�P���� D��rP�([��b�!+0��"�?D������L5�09�Ȏ^SĜѤ�?D��z����u���(���K�l?D��!w�P�,�B���Tp�D�֌"D�01ǡڂr-.ԑ��	G_�@1�+D��Q�jH+� #G˛	-¡��`5D��3#��I�RH-v���Qѭ4D�`rBJ'Z��v�ɇ۞ԙ��5D����Ȋ:ڜ��I��Q��%�#)2D��s�D up̀�s%
X˚}I 0D�`�a�N�H�lu����7�d��G.D���p˩0e�M�Q��^:B!k�(+D�,�6�%޼�:��ȿ%I
*D��g �2j�(`Ӆ�E�N�4ES�:D��"q�\�Q� �q�M�?dQʥH7D�؃���$��h�r�O�TZy��3D�����Q���v�[$�8���3D�T��ʌ�BQ9��&7�t(Vf1D�|����J96I!�dR,yrrĈQj/D��R�#��V 8Q�Z��f�2�-!D�|ڔ��*��U�dL6�4�c D��H$g�-i�<�iQ/9pQ�1�<D�BcO�$'!�Tm�(4W�@%	:D�0��g !��R�gS2�c�8D� ����	�Dg�~��ys5D�����;v}�q	��υDÚ���2D�`r�DS�S�K�0,U�32D�(���	<$��h�D�2l��S$�;D�  4i�m�r��5*�����.4D�|ۂ/Ecʾe�f	V�[��]J��1D�t�a\�i8��V�:J�	��b0D���D,cg���g7���pD*D�Ȼ� ��'�ҭ�F��YҐ �O&D��h��Nؐ�cA�J�2]�����#D��2-A��P���ܙ@A��C1 "D����)
:�(��Y�	�~��� D�<s��<@��$c��=Ty0��<T��� �ͣb]������@�b0�%"OJԹFx�N��#҄`�Ĝb�"Of��ڭf�����erR"O�}jQ�68�2���O�uF��r�"O|1	�fŌX���)cR��X�"OY������ <x�LB!c~���"O�0T�R[�q����4z��"O� �������^L7,��D\� �"O�E�!A,���x��~�y@"O69���jR�����ϞM�h��%"O�=���V���各A߰f��D��"O�uY��8dN��A&�d�H�"O`h��D��0�@�� ����"O$a̃�P�H]��oǢAߴ9"O�����Цc.��ط��4#��]2�"O��	s�+)�x&B�$�Z�"O�v�0\��-o0A`$�'OD!�D�V� ��/χ!��t�C�'�!�$Y��t@)��Fg>E�u�0�!�$�:y]r0�F��h���f�Wr!�D¯��D��G U�^}��k>c!�ďo�H�R��9J���Q�ˁ"�!��I��JUgW�;�� ��$�!�$�{�.̛D̖�l�&�#K$�!��hU�DY�f�j�8q�T�e�!�$F\.1�H�&~�B�&��u!�ɞ**~��@�y^��i4D�`!�� �pR���dK�.r�d���:zf!�$ͥ ?��+7/H�a�4s�ͦW!��y�����՚xX�V�Y2Q!�d̋"�8�b���a2Y��n"6S!�ѵ"��(0(^-fK�@;�J�+I!�DS���3�߄�h�R��B�oO!�DP�jl�[�+�4)F}�d�*Y!�$ڞ)�� ��2-p�С�K�p�!�D	8N2.�5�Ak����A�u�!�/[hB=! ���@k���4B�B�!򄊖qӼ��E�OX�KE/ 0{L!�B��+�i�S��eHv,�9!�d*뎍[t� 	�	ff�g!�F�T)�5��6,�~�dFɮ�!��(���r%�[��,�K��F)�!�+'a*ŋp��`���"r!�D�%8ɨ�q|�Ҍx���7!���4&%RiXq �;=ø���K!򄁶b&�����~��<Qq� �[!�DҩC@��a�ɛ�:���ʅTA!�$���E�Y�z��*Ri�mB!��&L(A�%+{a����V(��"O�(��M� �`p�dIצRa"ؘ�"Oҵ1���&w�� �56�ē"O4���ő�}���H@m$�X��"O�Q8�m�XXؠÌ�$Qi�"O�-�J�C�a���71pr�0�"O�2�h �x�c�ڂRh�t��"O�������C�\ Hz|��"ON��R�5jp�g�e[n�*�"O�5�d��4qb��2#ݼ%Vh[!"O�Y�``|������
/$�437"O�@ن��}bm�Oʹe"�8��"O��PJ�0��8���I6w�xA@"O-��*�gL��0����9"O.�"�s(L��F��J�}!D"O Ҥ��&� ��q@bܑ"ON��'F�+[���yVLa�C"O"�CEϳi���$J��T����"OR�J���932��t�6�j�a5"O΅����Cb�4HR�	~��"O��rV�ţV0�&D��(H"O(�x�[sƥS��^6a��� "O@ذFL��\��7J�^���[R"O� �5��)$�P���W�G:B�1�"O|�"b����j��X2��"O2l�A�W�aNdXx��	*@"�"O�(��Ȁ�x�TUzu�y����"O6̈2B�������YQ�W"O"Q��oْ6�A`�߯a�nQ"�"OАB�H+O��=k�_K��(��"O`M��R
i���H��.E��q{�"O��6���-�
`�S`K	[�h ��"OPԋE���L�r��/���5"OF=����%X�rAuKQ"�<CR"O���a�e�R�86�����"O��@ cόs��lse
F)V^V%�A"O��wm٬d7�;U
�RS�9�"O���@g['M����5B֑�"O�p# @�f������yX�X�"O�a�E�/2��5���R�v)v��&"O<�{V�W�vH�#`J,f.����"OΌ�%J�bx���CM�r˖���"O� G�5J2���T��"����"O���Kr�\������� �"O]���/����*����k�"O9� ��0�b5�5	C1��)�"Ot�e׈��	�h��2�"O֩ c�0*z�1Q�B�(at�k�"O��:w�B:�V�a���K,���6"O޵�!�ǅ-*��x �_z(��8�"Od�c*W������*̺! b�S"O*����+cuJ ҁ)X,'f�EsB"O8y�l�1� ��TH�4-�\=y�"OY q(^#f��He��/X�¬��"O��(1��f���S�+�4O͚	I�"O�Db���! x8���� q��L8S"O�x�ߚW�^�҃�[�O�ܥ��"O�Iɖ��<&�H�K=�R�� "O"����)[��!��QR�"O�a�W1	~��(�L�
����"O\� �����D�a+�4zJ`g"O�@��	�R��� jӠY��bd"ON<z�_���*�)��-$\�v"O���eG s/��d� +ya�"O�3�   �   !	  �  x     L(   �pA���D�Zv)C�'ll\�0BLz+��AI�o�'�|)��>9�D/m�$p��i[���=RU̘�_�D��*J���>)gl	[԰Lp��� O�PXy��(��!�Fo���>�f/��@�Z����ص?"Ĝ�T���&� ���ɟ8'���	͟h�>Ar'Z�p�L���]���P�!f�p���N>Y�ͅz�0 i����|�
YAo�zЉ�����u����  ��Ic*��Eņ�o�2$�ĉ�P�R2c�x�g�*�	M&T.h]!Q+D���1xsKA�L?!�RC��e �H��Xq���g#azr�d��\��)�� �E��tP�
!��?z����f�Qk�9	҄%��O��EzʟLT�BN:k7�0k��)H~0��wd!�=U|kd���4��96p�,)���,��<� �xZ1O0P� *S)����y�h@��ӰuI�؁1����ȓm�V��'�V?��qI��������<i���)]�5�x�3�Vq¼x��]&'b!�D�	t�� �2.�����[�	�U�"=�*��Q�?��(��g8��W �6~�N8�"�՟dz�i\"��'��dF�����s϶�֜�� ��U�l�Е
>��?����1B.uFeS��H�@�PH�<�E&�==8H	Q�\$PC�d5ay�'F�y�c@�i�T�B+�CG�� g�&�y��וx��S����Ib⩩����?	�\����d2�	*9 �j2͒�e�ۖkY�m\��Z�l�������p~�L[�j�ŋ@��	���P�o��Lar�\�� ��u��rGa\q����g��}�e���6M4By��L5e���͜;ڮ�9�E\�At����\�����Ly�'�O �$��22p(���E6 8uʱ�'��O�<(E N�x�h�a�� \략���ߑK���d!�i�I�"D�(1��
.[2�P����Ay1�ȷ�' ��O~���ǳ$n�AAC&4�|��0��e�<�Q�PJ1�B9%d@q�FGnń�	u�?�F�3r���N�B愑*k� =�����z�ז^B��QG��@�m�?���)d�ߦ@�����1t�*������'N��R F�C���S�O8Th�lX>Mn�*�	���l�Z4�>��.���� ���T�D�O�����L�,Qz6
����'�,�;���)�"_�D�{���t�tUM��'(�����?M~N|b6�W�'o̡�E�P(3�`C�(_~��?��RR�8)�� .���K���	2��Љ�D�?�ã"(���a��������t�4�B"j�;T¾�l	[]��:G���M���ަQ�)	r�D�|:��a΁��7-u��N"1Jayr(�6<=���K]$<���j��ؐ��'���˓`�б ���3>��BI
��0�*=��Il���L<&#`����H�2��(q�!򤕜afH�1!�=
��#�R�u�$+d�2��?Y2L<���k�������N�	��l��A�p�`u�q�����O"�d�<Y�m	��?��A��$�!�+�li"II�O��P;�-��*޺p��I����#p�"
�e@4nɧ/�l��NV#0�d��Qhr�F�􄑘m�f4p!��h!�������Q�'�R�8���O���&��=c�*�Q㛾Q�B������>ɱD�v}H/�IA�ePMP��M)n8�ypo�17s|&�� i�ßh�'��5{b�1�I��mÀ	 [sN}�t�;7V"��#Hζ�?1-O�dKpL�O���iq��[$��i��"8��B����ȕ����^h��	�#x �t�W�.O���V��q�b�M��c�9 	��I�:#�$��u	�4�Mu�1w�B"�
.M�nu1IQ��I՟L�?��d�;pRPcR���X��{�M�S�W���4i����%���F�&av��Ŏ����'r�As��45s�'����M�۴ψ������"5ӥ$�.��2#�'{�l�(l;�%�w�פ������O���B��{Yx4�5l��=�b5���x��U�[
]kGD܏b=*;gi%§q�𵣒��`f�Q蒹F��%��*���O�DZ�S`�)l�e��U���\�� 3'(�����UX��,1�\�Xwk���J��m]��ۉ�ϓj�R����i��'�6��3���WH!s@9)���;@�i0���Igy�exG�7�$�S�? P��bG³�l<˖&P\��x���01�T�'�h�0��VQ�$B�7w�բC�ܨDҔ�Q�ˢ�'H(X�/�3��H�����7���Buᔴ`�p���t��*U��)�<q�4�\�ش&��@������ Q@�O\�j c[ ��|��%O��ˡ�'��	8E� "<���?	�OD�p�j�&[��AA�C�#4z��O:@mڻn�ģ<y5+0�ė3w ��!ӧ4�bո�`B5�!�ϴ	�<��Ԃ�4)��e�
��!�N�J^�"۸\����.��^��C�I1|Ⱄ p*J�os֐:BEZ�ps���
n��W�(�)�
"r�yQ����8�G{Zw� �C��%!���i�i�Lq�
6N��d�>�3E"扗'������8cm� ?����Ц�[���c"O`�+�,�0O���`O�:�|��7�'��O4����a0l�@&N�`pB2"O,ڵB�/.��i�C�#��f���S����Ć����L!@�zq`�m�'Y�laɈ�d�Wɤ�<afno>����k��%:D��7`-n5��)H̓3tJY�b�=�3�DS3�D4[��+VL^�a����~�!��Y�*���B�Y�\H�H��bS/�1Ob�=�|���@4	�8���H�iU��
�p�<��E�jv0٩ac��g�U�@N$�HO0˧:��Om:�U�g["�H��Ǭt�,�AB�'Z�A�-�I'Q>�d��4+sr�y�hO�Amd�F�<�Oک�pA-��][Ơ^
y2�"O�ɚc�XM��i5;,hH5���Wx��3�+[�zr��-M�	���1�A7D�਑#E	�z��t/4M�n-P@��O"��'�#=��yg�c=���;;~D���~�B�tAF�MD�'�r�ʣ˜�3�Bm
�AΫ4P��
�'sL�S �3G�:0rԌW�A����
�'�2��R��)��H��G�5=֕X�OR�ʶ�B]���@�\+��9c�'I�OR��U�� (I�� 2k˩Wa�qW��"�Ӻ�A���tA�L�{����`͉j�,��7N'��;�1O�!IP��� S9�.b� �J,��R����y"
Da'��T��̊�L�0=)�"��^*%�1EPL�������yRS� 4	"�:P�ii��S��'g�#=�O�ƀ��V�@Ԋ�(D��:Y�L��ɧ1_>�H�y�/��|2XHc�uJ��Ք3�L�f✈ј':��g��n�g�I��Ti��K,? B :A*�iU�C�I�yy8�Qǔ�����
T,��b��G{���F��R�hi+'�¨4th
�`��y�/�-����C's�RPc����#(���OBr㟨+���u��y��UZ(p��O��p�o���|�I�{i�01"�N�;t�<`!E�\-���G�i��x ����pbQ��vrV4C��,D��I��P���H%	���9�.���<Y�уSٔ]�2	��W�y�Bl�U�<��kM�$'�݂`��<�d	�fMӟ��O�lDz"�DϠ���P�� 2\(�G�s7���Ѧ�[�,:�(]�O��&烾*@BLJ�Ȝb�!�"Od1���l�R�;O��YG"OJ06�лj¤i�2+H�%�\j�!"4�T  hֻ`�h����I%5~LqF�=|O��&���EM�;[��e�ȭ5�ܬ��'�I@��uW(�0�?!�GR�
�dr���JQ���D�r�q�zc�t
Ai;�iR:	m�U�����v8� �=Y�!�O��I�胺zr���ꑖ(�az��d� 5p����㘶& 4c"*F��!򤗯B�^�T�#2����"��7�O28Fzʟ*�3�¨#�v�2�	�0fU:��`)7ړn�r�S��Ů��$(_�n�ZŚ�ȓ�z�"`���I*�1O������
����S�? �I+2��d
�aP��O1OJ��K�"Or��P�I�e4���,��*�P�KQ��5�S�'r���#��� T�g �gQB���^O�ѨP��2o��ءV�$@1��ڌ�d�|z���*%��L��jҬ��{`ǁ^��@	� P�b�X����OFСSd��bux&2f�yA��t�r���@h���9TgM�W���`e��-#!���<Ŏ��鍟sK�tA��W�����	�9ð�����Z
��`%gc�C�(
H\���,Cx��� :NK��$BW}"�/ғ��'�M�3F�!�^`��Q�H�h�'�B7�)^Q�8S��|FǜZ[�j�b�X�`j��)�yba�|��D�Y�JX�	t�Y)�yRf�4��lB��� ^%�itO�Eӣ�ʯy��H sh�GA�$(f�'���Ot��S�E}��('�F�o涁:���&�Ӻ���@��0ş?�J��A^5>�ـj=��4�1O̩b"���iC����vM��ؐ8p��y�-ږ(�@�Hpƾ �D��G�0=y�B�
�^�s�δ�(qǀM�yR��[�"q�tܴM�F�# ����'�"=�O������\�Z��5/�cR���b�	*�����'Mx��'.����1)^p(��b����-��y��וD��M�}&���&ɇ���*�$r\8��-D��h���Psߎ'|Q��B9�l���OZ�u%��ka�wF��O����'.h��n��"�~�R�7P�: Ѐ�k��E-�	�d�� $�ީHH uk.
�8�J�?�`�<i�*�� 
'ބ)�y�Ue��p@��6/^�@~���	-1��� �U1��rP`�M�B�q5c6	^0'Pl�9�
�H�"<��+�%���o���w*��J[�Ņ����Ń����`�?P�n�������I�'�1Oʐ�$(��"��/���j��O<pnڔ]���<1�o1�$��i���*ei�<0��vn�>!��W�d0��mM�x6U���u�!���D��*V�_}� ���S)2�C�2U1�x�r��`���V������G��)��H��O?/M��m����@E{Zw�
����=��	���.��@1j����A�>��(>�	#,\Β���`�H#���x���1�h|�"OFP2 ���R� ��1��;}��؁�'s�OI�WHɨ\��u;a�F��.��c"O ��G�艩V��+?����U�$k���iF*�.���	�t}���2��
�l�=�b�4�1OF��O���2N���D0!��:���q� t��m���L>����4=��ۂg,p�'�Q�<)��	 b���k�
�#wi�-�6�f��hO1�pA16a�n��5��EZ?Q��#"O��q�i�KּD$_&a<.M��=ғ���S��Z�GF�6=ʸ%$�
��Ɋp��(�yrc�J��?�V'ʋx�鉶�<J�j�`A@P�Iu�P��0�y��e�F��VO��"��!��q\�=�"��/ӎ�H�(J>[���Dxb�'��Ċ�I�/��,�P�L�m�����'�Լ���:i�d���Tfk� ��Ks�I.�HOxc�����0v4p�H���`؂e��|xٴh�~�EyrJTJ��	}��횉s|n*@�ڶ]FC�	�����V�.1���[�;��B��<D�X�+B��>=5�ba�6Oc~��Ɠ=,�zb*_�~���q"��=,J���I���[�U�%�@���1�䂠`�F9�?)����Jp���''z���H�33N��D
o��k�}���q�hh�'?�r�Q�2�Ђ0-L�5��р��0D�� ���D/R�e��Ey���Jը�ӳ�'�OH�*�CHu�ؐ��눒` �J "O����,�)T@�6E�U#��dQp����GoRDb��P!l����u��+�(�=!� <kn1O�!�O����mպ֨};��P�jI&�$ӝJ�`��L>�@%7D� 5�6K Ph�w�<�`�R`H���2Qe
}{Fm�u̓�hO1�D��eԷGaD��J�!�>|R�"O��J��@9	7Q��)�،dY��(ғ����]��,PL�A�}�t(ʢ�C6��)�	�ˮ|!�ymR��?��&���\ �c��<�p#�j%o�18�t��8��åf
��Z.�YEȵ��Zܙ�4d��  �� ���lܤhDx��'�H	����H�U/ȱSI�q�'�(�q�P���`����+�9��x"��<�HO�c��
[�X`� Eň�M92�����0��4/�r�Gy%
v�ɵEgJ�2������ާ<��C�	W0|�Iӄ�=0
�H��]7�B�I�"ز�`�B8�\@�Z�Ndv���u�]U��j�����˶^�Ľ���"��w8���v���N���h��>`���?����>���'p�
�^)y�ȝ��[���C�}��d̓1$��&?��S���V�@�P&ܾP�7+D�����np��q�
WEx&��Pn>LO�H��P-?��\����:4�Ap��;D� Z�����M;wl�{+n��#;�I�HO�S�^;�8"1hK"��)EC-� tE{���Tq�c��a�=�((�BF�?Quըac�AҪT*�+0�k|�T����|��D�o�� �A�M���b3ė��y��.,�>u8ǿP�!��4�$���y��)�3	��13(�T�0���#�..�C�I"I�����D�`�^(S4,8EzV>�)�"F�u�°Ht�
,n=2���?����4;�1O�a����'�H��sA;'::���.�kf�� [�B*�#��C`N�y�>�ժ��ybk3S\�� �bI.pc:�0�e[��OD��d������Xz(���ҋ!�dm�8\�AdG�_\j�R��ߥ7�R��>�1�	W̓6@|�@dIY�w��A�+8I����-��� ��(OJ>�u�F1.�)b�[6� ]���Er�<y�E�=5T��Q�	/��صhl�<ᡭV�H���U6n64
r
�'��x���%<Ը���¶��HI'��7��=醞|��B���(t&U�R2�S$�$��'�ў֝�7�,�䎳v>$��kY
�t��3C�O���y�g�"��'�R-qw'ѥ"��R�T,e��'X���S��- \�� �ɗT�9ӓ��'&D���������#S�2���'#�P��'H�O��h�jّ	�v��B9�S����<xb,�� }ϴ�y��P�ўh"���!�'�h�'b����$3vH!���/`�Ny��y҄D�r��}&����&u:�Y'��b��h�..D��IC�3��<�CkQ?Be�����*�Iq���O}
���@ uY�GԱDk���'�J���yD
�AZ�f���������%�ɭ`&���u�C~��X��� ����Y/%����<��9�矼��CslzI�6^e^)���?.��	����q��҄G�*U"g@�s#�C�	�tڦ%�W'C�g�.DЕ��2�"<iϓeK��d�ђ����;��A����-��}YZԣ#H����	����Z�'�1Ob�Y�FS�;<9)5�҄ ���kC�O�mZ,-�Ң<Q5�4����qVzlR�P�`��-s�KA�
�!�D�����pv�N��|�/�35f!�� ���J��6��@)O�M�l,ZE)4�X�P!�=����["��i�	'|O��'��2&Gѓx��R�ګ�j�*��7�Ip��u�)P�?�#Q�a6�d�T&��s���BC�v�5�c�ܓ��3�ɔ[tB�!�]�#�n�a�C��E�!��B�[`�`��n�F�<��!�h�azB��N<S���Gnș9���!���!�N���]x���� y������(�S�d)4hBr D��ed\�Y�ܼ[eў@���E/��'��Aϧ��hI6.�>WԦ�VM��EP�K�yR���E2��}&��S�.Ҩ6,�`s(��xB��Za�3D���� ��\:�1�'�d���%�,�IE���O|H�K�/M4@W*�lF�)1�' "���2YF���.E�h��<ە�Z��!��5�|IV!E�(9:��b��y>:	����H�IП�����M#��?�����ĕ�L���As��$��E���sL� ��؅+d�r�� ����1����sp�didޏf�ޱ�c&�29z�1�D�%$M!��O���&JF�g�	�\'�cG���]^�8V���J`Z���DN)#�O����ȃ]}�����3Mg�(� �1�!��&,	�aӱ ��H����5���l���C!��?)�������C 1����dBD�$�µ���u#؁�M�Dn�w�'�0ХO�a!tP���s����BɃ�mP?x��m(�f�������8<O~���Ԅ%��u���,%�PxcR�8D���Y�,W/I4Z}��)<O���Ҩ`hb	��ό�g켁ďI�C���'�ў0�>ag ��Vo���
��N�P1���o����O>�bܵ4H�8�@V�fE�u��_`�]�ux����]�%�p�Oy���šP��T9T�äX������]#:l�Ĩ<��?q�O����VXG P�4�b���������Z�J�Ă��+,O��C�G��������<)@�� �� ʓ�Ӱl����cIX�Y��O����>��U%ky�x:��_.�2��Y~�°=��ƯES|�둎��QB���I�A��]瑞�'
�lI:��(�4d���@�i3�ܘUk�$�?�(O����V-����'T�S�M��4(.P�I�hL$���.�}VR����'�ҡA� �^�C��_�]ԧ�ŀ+��A�Ӏ[eH�8��N?����s!A�4��O���Dϙ( �sbmAq�O[ �A�#J�����Q� �H<�k�����IO�O	�	^nX�	`a�W8Ds��yB��_Kb��#NN�:t;p����'g�x��?I�K`�(���E�BFpu�@o�ڟ�d�#D�'��6����O�[��>aUP2I)�[��yR�����}�:��d�e~e'o�?v�!�dO�,�h�Бn���!˓Cھ��L��ɘB5f�P��P��A[��6@�C䉶cD	رx��p���q�T�$Vc}�I#ғ��'C�0�w%ɮ(Dx��� ̰^�pD��''>6m�$�Q�̠��|b�ա=�p�v�H�r���!�#A��y�B�6Kʬ��ҧo[��XDˌ�y���.~�0"��R���	�d��?��B#B�P
s �%D�$�hM.	_�{�#$�$5V%�E1�ҔdE�=#�E�XB�O.�=�;1Nzy�Iq��UPFe�;9�FQ���&�c���{%�
��!K��1�M����CUm�0�@$�ȓi{���J��h&�<*�M�k��IS�c�<��g,:q\ѹ�A�*l�q�ȓ��l	��ɿ@���Qp�#o��P�?a���?m����0^O��Q�"�P��ѡ�H~�'�l�H�c(�ɡ&��/qTD:fM9Dx(j�Q8u\�b�`[�&T8.�q��'>����]� �����$ԧ}���'Wt������Ve����E�	,V�q�y��)� �.�G��&	�]k��8&ʬC䉿à�c��<��qU �(D� DzR[> ���!}�����7o�<p�GOA�yR�'m���� �����?A�>   �1��A%kp��.ʆJ���*S�+��y�h=�U�Ld�y�#�ce�@̓^��1��ҟ���'���
&�*Qyc)�;/�h���`��&�!�$ׂ)��ٳ�썆JR��B���+�qO�ϓ F�Dx�'�&�R6��l�+��	Iu�'%�'V���%O!)���'�b�'E�6�+e��P�r Y)<Z���5�#b��9d˞���D�#�Ʃ��ĩ}��3�E�2�"%�E8"'���D^�Q�� �\�P@�C��$#�K,Fx"ė�i���AńI��晒��5��d�6�'Jў0�;t=�a�_�qLptnq��oY(<�F�	�,��ـ�H�6{�F��$�U�P�z��A2(n����쟰�<����$	���0 ���������'W��i��%扴}d^�qUc-�I�:���ƮP��|����?Vzԑ�G�<�w��S%8�Q�o^�w(�郭�E؟L��}N��ǧ,N�Xp�R�P�\r����i��X��������t�㉞�(O�u/�±�dHʶd����#�(��%ʑ��c�'Ǉ��p�$Y�L�mY�K�s��G��Ĩ#���P�e.>��,z�-�� �O�0d�{�<y�FQ�$!D�"8D�4&�x�'�Q?ň0��/>O6�鄩�
����:D�p�c��{�E��)��	'�e�S7}��/�S����X�1Dݎ/�
�� �?3�찴+3�I�D���!�y��'���I�<��S�� U���W�Sp��ʓ$o�<P��b���q�)�$N����b�0%O=D�<�7�
�eǂX���##��KBĹ>����3� �XqTnJ��}��G�&dJ����"O�1ʀ	R�pi��А��?gT����l}BD4�F�0��E�?�H���J//T��(�h��'�1O(P{�%�w8V� S���zԾ��kV�Y�\(ŧE/HR�e��5���J�*�$S5��W�C3)΢���jX.� ��I�+
$�������9$�4��ɾ_���]�(l�@��F�B�	U����a�?I�`P���"�^@bS�OބGz�/� "� `k�Oj���o� c�*U�ܴj��0�<y�G��j�t�<� D��j[��؄�9]�|uӔ��9�n ��'�V1��`0`٨� ^^�������~����fD��1ŀѷ;,�d���y2$K�\X��V��7�@r�/�p<A�創m��}�'h�-o�T�� 2�j�'�hb�@���\�[�,�I���ͧr�,�lյ)隸��d5N���'��5zЈ�Oh��(4��p@�����?Z�FI�pX60�S��2ڠ�r�j�r�'l�����W�)��cH+t�h��@Y#7���J��"�� |�t��0BDu�T�����ȓ	��i�u:(��Q�S?���O�AGz��|`��O@\��PyK���ֱv���P�(�	��ZM>�O���H��O���VR�>���S��O��y+C�Y8��I� k�irLhS�޾l� xD�Q(%��<±䟨���1�_,cR�i����Sؼ\@D��!E�D1�i�~�Yw�h���a?�Zsf�#�S
����ŖuS����M{ �[K*ҧ�9O�p�AkN�; �P󈂼x�$��H�vʀ�x������<Ab��w�d���y`�֟D%��(X�x44C��yaK���0�Ojm<AMB�}�B
`Yqv	�7���X�	�c����� Vj��S����3O�E��>��GH?N<���ۭ	#�!!oȃ����dʟ̢0/}�IG$!��D�t+�/m�Y�C�H��r�Y�*d٩�N�5��I1�M�s��J3�-}@j�x�r0
��O`Q�Y�/0�}* ����yR�@���I��M��.�'Q`t�`@�·-�JЛ �GN9�H�is��� Œv�T>�ɽC|��@]Qď_g[�ݻq�����b)tӶ(9�'5��A�OYi�4J.�>�	�!1���b`g�(@�q�g��O(J�4��E(?��y�lھ�~�M�'��9�a�>�4�	�?Q)}Ӫ��32x82�+�� ^��+�B�kld��4`n��e-� �^P{��͔D,�n���%�x⭟��Z�ܴu�Zdi@���Z@�1hUt�6��'�'��	G�	f?�/��1�*��D��'�	�@��Q�<a�!����Q���1uhѠtXP�<��#eԜ�#�x��`AiHN�<�1�i����dH�A#�1���S�<�`��{q,���h��X���D�<��� 0����Ώ��J�
� Iz�<� ��S�bu;�M�5PY����n�L�<�eX-=(�	3�Ӫl�NMq`�DF�<	��/Z��0�f፣L0b�1�fRI�<!��Ę ��|��o��[)��	g�\]�<�'
�2�tT��jV�a�$ ME�'P��'"�'lrPe~�Ej�	F-�X�ȶR��7��OB�D�O��d�O���On���O���/T�̜��ѣtU"���ŉG�v�oZ۟d��埬�	��@����	ğ���b����2i�y"DE�
`�5I�4�?q���?���?����?!���?��,���"�@�~�����_�4+
�ԴiP��'�r�'���'�r�'���'*��a̕�W�4ѳ���,v�N���iӚ�d�O8���O��O��$�O>�D�O�R
�3���g�" ð�sƇ䦁���0�I���I����I쟘�	��hs��Y4�ٰ.9E�01�����M���?��?���?y���?����?)7��^4��iFŗS�"52T��f7�f�'�B�'���'�r�'���'���f���o��- Yq��؆07��Od�D�O���Ov�d�O��D�O���׻H0� bEKT l1Kâ¬8ml��|�I�@�����	؟0��ʟ����G�R�#�+|����E&{j���4�?Y���?����?���?����?!�Kj2h;�M
���ug&sI���0ƚݦ1��ǟ0�I؟��I̟��I�h�	���F��5A�h䨧-�StI����M��'��p��#;���`�4�D���Y��=���9%A}�c4,�ի ��0��'���I.������λK2��բF4**z]B��<-ڐ�I۟���%�?�U�ZB���h����ZwT��'�E�#��Ia%�p��J��P�V���3���	�$���Z�X���($���yBm�9e��-����,�P�h��?Y.O �O��q�@�$H1O�� :��j����j���
`8�'[)3�O�=�'�'���&��O�8˳�Cv�zs���D�ct
]�X~&8�'{N6m�u�x���}哽EE��$��x��s�P�[�P	�'-_� U�%�9��d�O��Y�J��;(ʓ��d7?) '	$��!��4A���h�ʟ`s�A d����'�UJ�����6Qw8<#��3�>�x!�ߩ|
�Q�(��x��;p�,��g��1�'q�t;�4Q�L��m�n@���Z�� `X�n��<�5M"gc�I�<�ao�����9.O��'h�d{�H��tAp4�pᛰ<�.�A��	|yB�
*0z�}y�y��Ot�i	�O �kW*�=��}S�gc��I�V�y}��'��Mʎ����:f@� ȟ.]���<GM�M�b	��.��YU��"n�{/�~�h�*MW-��# R��/O��'�p�N�}}�Eqvh���>�C�Z1�8=��'�r�'L��'L剫j��ڑ��$�c�O�d���F 0��1���۟�޴�?���a~�!�>�R�i�z7M��f�6L��8
�\�p*O�I�蚓�ہ:X\�x� �?��Ҥ(����T��F�~1h��]>a:�w�m��56H(���N-k�80�59����?q��R��E��'�?�Ӈ�%�,�����
E�;17�?q���?��@݂&9�����?�a�i\����~��V	���0 ŏ_���b�ՑS�V\��t����G�Ï�M+��&�)�Xw=
bT!RGB����4[����Fh �E�G�a�
-�㍓^,��1Q�,�u�'8>��[^�98���?��&��������9[���D%���?)O�8�nP�,=��D�ON���bm�� �n�Դs�^8(P��a�E+���iG�	��n�wf�	[�BY�bߟ�(��"p)�V_�+��p�󬂡r�|C�	@��M��Z?�G	�Y�
扗L�B�͓��&�>Q�T!�동Z��4	2��?	�&^&)r��?���?���򤒉GX5Y�T H�D�T�IW�4�Y�=�Ԏ�O��D���e�	�Pg�r��	�M#��W�2��
 8hU�AEoT
��J�Q��٢�V�u�4ͫ�'�B�e"U��o� ��̓T4P�VG��.0��2��!h>�P��?��o�2/�DXJ��?Q��:�E���)�:<.)!�)M(z�v�J`I�WC�0%K�~����S$�"��@�4�y'+&L�R��Ȉ�}�jh�S�����y�r5��O����������.>ם=8�4��$z^��2��S}����GIV��?�wF�>�6�I�Y�B��{6`����V�:�5�����Z�|�F�j��C!f��;�"D
!�$�O~�d�O
�h���Pubͭ�?	���?�t
ά9}p!p&���>@r�এ���?yp��v~��>yb�i�6�L����t��jr#�3`��Y��ͶG�Е��N"�y����i����i�8�0O-� LN��y� ȚCvn�b��"z�v����R
ה�ac�O��$�O�$Ӱ^�k�j����D�O �	/1����� m�r@ʖ ���	t��;1��O����]�I �Z����b?6*���E��24��a�DC��a`���U�vFu�n,p"�����(f���E�#�i4H��'{������]�� !�M�Y��d�j�����U�ؘ����O����O�����6q��sC-qܬqѬ�dID�HvF�<�� ^�1p0\2���?����q���|2��e۶'!xD@5`Z����Z����4�v��4�~�얈H�2��O�� ��φ"m�Q�)L�(q�����A���ƢI?���N�1�0 �'{t�S;O� ,)�(L�	@�0�՞�~1����>�	���"�'K�'�bY��e��J���I%5���"�	E�k�d�j��ͺ�%�I%�M[��m�lh�'����?ٴh4�������A���&Y��a�E(m	�iPI�'|���ϓ\j
p	�t�7m�+�@牯BAF��;o�@SJL�:"�Dh����Z�Z�Pp�X�!�j`�	͟��	�?�`��Q�S��P��7��h��[	f��xp���t�Iɟ�b��(�(�'�6�O�Y3��O�$�'b�!`����IIpo�|��I̡�~�cSg�b�y��i��Ԇ#L��NX�f���ӎ&�v�Jvn÷s9,YeJ,2�[��R*�y��"O��$P�5s&����9�a�!�OT��O`���)��:�2��T'�r��O���<i�L	�A�B���?A���2��A��	Jpc��P�Xԯ��A���)Ox��'�7-�-�ᨹ��s�ėnA��N�Q���CD+s���1fV�?Bd�`{l�� @�{bYȱ�NP 1�W���Υ>�1%�a�0b�}��P�p	�X�$l��,K��1�-B�?���?���?I(Oʼ��Ju\87I�>N����GȒ�Pg��<IӺi��b����i}�F|ӈ�1Wc�H�"�(Qh7~�T��ӊBܦ���A+/_�I�"�����0@Nz���FJ�y򬍎%�B݂ψ�.- ��	Ħ'p�蠕�'?��B
'���'���O7ґ�W�?q��44��(��-�1J`ꈻ��G�@k@�Ue�O �$�O��i�C[�ʓ)�f7�0L�gD.��(�I	�Mc�ɑs!c�p�l��F���	I�0��^��)���ؠ�-i���ʜ1<<\Y���+�*�S.Q02��3��2���O$[���<I3���?Q3�*$��� �r�A�����\��gٟ��j��?i��?�(O:���_�\���O��D�5oL�$��EV'���3�(f��,��I��J즹a۴&����9{��UJ6af�zec�'^������牯sf� UL�9�ةc�y��re��P������e��ߠ rx,{��]��0E`��\ܟ�����Đ����h%?a�Iğ�͓@6� 2�I�?)L��7�
?��H�	2F)�6A�����%�	x���JFoT�p�����t%��R5��	$zZC �I�ɛ��Ĉfi2��A��t����h���4��/9��^*t�]� @.��|��D OoRQ!� �y"��7$����&FQr�!�'���'E��W%�=��R&#�h�k&/_��cAT�|���E�]x|u��П�I�?y�eg�Wy�&��jYu��L[$�@��0�˓�?��4,�<���2����7&2��>:�v5"5N�̄����Q��s�,��V�̓|� Ő�m�Ov����Y�<�'���?���4y�an� U{薋V �����?Q���?���?9)O�-Kc�X�d3��d$� ����]*Dt�\{m@.K��Q��'��7-�O�42���C/O�D~�����`������"��+*���D_��%�VmJ����X�:ONdq���.�uקF�	X��Γ|��w}�,�d�̝_�RMq5�R�z�m9  Jĸ	��?Y��ReƏ��'�?���<������rr^xʴ��?a��?	���L�e�)Ox�oZ�$�Q箟d���ēOP��EB�L���:$���H���ƌ]�A	��w�.�I�6A�ݕ(��P̓
�L%��*юk�2����A 9Lĝ�����d�4�I�m��M�	=��H7ob�'�V#J�Tk�M�y�a�[�E�r�'��	IY�pӆN�������$�S�!b�p���=d�-P@ _��A�yy��>qE�if7-DB�d$!�(-A�O�
0�U�>z��{��y�|	2�
�R)�P"�,� �Γ&�
̙���OP
 (��<���U`�}�<-q���W��l���O6��E� wh����O����O<���<�ԏK�u��H�	�1x�)�@�\��i0�C��?	������'��T��O2P�'y��P�Y0 Ƭ��pۆ�P��ݤs��%�/>�4A�����^4a�'Y���S����oZ�y~�h��`8,xi�/߼j<�����$S�HDnZ:�?���6�@U���?y����!�[���)àF��q뎅(��[�b�\7��{�b�98���'%��O��1�O� x��杈j����4�	mU�����b ����O�����O(��5-����IB�N��C�rP��;b-FYBh@��ZE���?1��.(����q�|��'E��dG�[��m��O��w�F5YHܪ��M'I�u��OL���O����<y�*Lf������?���_��Q'0g�l��G4�"�x��h���'N`듸?�o`���HH�p�O�P��I��%=tٱ��/�<�	�Ď �@PѦ�����K�����y���C[ X�L$�0����K�IvV�B���O��d�O1��bVԒ�L�d�O�扛Be��$��m�~� ��>�*��4+U�T��<�E�i�����$�����pD�!�㔃>�R�y`��k*�@���O�9X���q@��VPUp��P_6)�Ga������F����Ћ�=�(���|�0j4Z�<���9 Q2����?����?��''Ί�{�K�r.�AK���aAK��(g|ɔ'`vu��͸D2�'��O���dT����D��`2+�h��L*������$�O���R�K8�DF�!��UP͟�\P2+%n�(<���� ij�(f��<n�Q�&�^�p0�䖢JI���n��Y5T��
��31�L����F�]���7U��1�TE��E{,Y���?���?����򄟲��ː��O��ݶn]�3JT8Y�-@fn�O�Eo�ݟ0y@�6?�]����ݟ��8i�03M�w�&��-�6K'�}H�̃�V����ʟ��s'��5���5TT3�'��·�À�:&p�Z� � #����@#|�h�[�����$��ퟐ�ӯ"�2P&?I����TiѰ��R��lrǭ"$�P�I֟ �	6R�,t�F�ПD�ɴ�M���x/�-~@�X�
�s�$2�P�&gڡ���`?�S"�+H���I�?���Nк�	�5r��)R����o�#���s�ibq( .���y�&�C����?q�E2d������?A�gT������N���JӜ"�����?I-O�P-�G�����O(���� a.yV���E�J�l��t����8��Iǟ��	�B���9aØ�du��^|����=(�!@���E��/m�|����9u�d��u7dټ�?���u'U��r����$bgDY�2_��С���?�4�A�{?f�{���?i��?a����@��6�a���{���R��V�=z7�ڏ��ʓ*����';����O��'��n�7::�K�-7Ğ�h��r"⃉�Dzځ��/�4�?��'<f�ID��캋�탸<!���5R�P�0"j���Fm�Z�$�7�˟\Ў��J��	����?%���d��nV�?!�D�A��5>8 1BV%s��i���	��?i���?A��O^\�Χ�?1��i���,5��㘁o`���C�E�4.6����0岟q��3G��*r@p��;������7�x[F��X�xEI�	ȭ
a�8�ɶQ�����>OP����s}�i�O�-A��߭U����ݯ>v%KVh��"����a/#6�d�O.���O��e�B��S��?����?��I���#�fO�A�q[��?�S��<y��o�����M��i���X�=O^`9'�E.p���9v��4%�_��'t@h ��Dh�T�f֋��i����	Tƹ��� �V|II�Jz�E!e��ɟL��џ�b7@��"$?i�Iԟ��.� �q��#$ti���^�V���I<�蓡Ffy��`��dE�hu�	�?%0�R#K��h��á�:�!\.e��4����� [�G�)	f\��sͨ���'�������3A�N��u8YH�sq���;�ȡ,�l���+�<E�'�()(bJؠmK��'���O�t�a�"�����ώ���	j�a�?M��,8��rOƟ��������'Ҹ���dj���>���g̣k�.|���Ͼ��$�O����&_.��H3~�v9X@�'��d"��H����U,
2R��|#"(\�I>�t�$�i���9O %��fD�yr��y��ɤ�?����JSL|�F2v��ҲD^�Ƭ�W�S*�?����?���?Q/ODДD��HH��]5MW��`S�FU�
LC��"&�$��Ϧ���26�s4�ǟ$nZ$j/������%da��{���=+���J�U?�B኉�Sֹ�I%W}ą����-=9��r�u؛w�R\2��ԘK!��S��l�0$؛�2� &���Iޟ�S�/w��'?A��	I����ǂ^�JKBl�`!h����	ɟd��%��H�. Hy��s�$�D-���V��vYA�ߨ8�¼� ˜`l��W8O2�$��0R�7-�h�sg�	�e��<�e��S̰1s�OW�y��̐'n � \������OF����DyrI�O�5��i� 11O8j�ϒ�L9�\`�"]:^&V�{3�,��W������I����ӒQ�Y�`�J�W�a��!��}2�2Q�Py�G�>)���?y��z?��倴8m���1�4(`�Ae��鐎�=^�1�Q�f�7-:��韠X�<O,��L�<yE���^`�fC�J0�`BeO�2\���;5cp+�'���'%b�'e剬{\��� rM���B�/PԜ��+�����"��/Y��'��7��Oz�#;O���V~}��'�1	գ�0T �	�N �b�'���
�9���6M�����jM4���%ٓ
L�<���\L�F��>{ؕʱ��5�M�w�'Z���g�hb�'��OV�]�P�?%�'�ֈ44�2 .�,d�	�� b�+�O����O��i &n�4�
{��5�:A�c��HJƙH��-$y�W�'v�d���~RUsxmr��Z4e�uHQ^
,X�`�?���0�g�($��d�O�E���ب�?!V�B*;D�	�?A!�!
�� ��bR��2-I�v����f���r��ݟp�	���iyRAS�,,�|�b�'���'V�uA��V�����[��cv�'�0���O8�'6��'S���'�* �Ӟ<~�zp�c7�dj��F"͓�hș�Ō(�M;�KP#���.c��<O�<��h�>,VܛTl�j�:Y�R�t����X��#�5���'?���şd�"V�"�`3�Ѐ0ӊ��c���	;7^x�A�ɟ����Ms�Ug���'`��.��B%0Tc�8[�f�����Y����"�,'��OF*>�:��б�SNl���׎�+�i��Yp��9^��1���E���IPA�74�7�?y�MV����q��?����Jaԭy��$�*��o @����ƽ[��ܡ)O,��IǼif���O�d���\Ç�<!�AN�!,��b�U�_�|�rP/�	�|�	l����W�\a�b�?�k1A�&�h1	���q��3s��?7���n�	r����1C�֐kc;O���➟P:��,�ެ`��ҙ:�fXh���"'�dsA��1Y�������?)��?�����EY5i��r�h��EĳQ` ����5	H�1�Ԧ�O(oZ�L�$�9?��\�L��4���HS 3�e�0i�8E��%��S��� ���,մ�BՁ���y@�PZ�}�;-�1��H�|��7�*<A"����X���ֱ:��+��s��Q��'O��'��&2D��OZ2g׬� ��ԓ`M$P����bLb�'12 /D��Y��T�`�4�?�A�h?�'�Us�^C�!9�M���{]��͓7��<�j�$�M�'W��t1\w�θ�'frj�e�2P m��T�[U���'d-M���'��`I�<��'��d���Hu��'p"�U�I��ف���1G��ˀ��I��'��I�
�ޕ
f㟨��՟���!1N�8jǩY�`�쬛b�\��a��vy�,�>1�i�7�@�%���	�}�j	yޟC������$��	0xt�p�ȵT�Ji� �X'g�*��'����<SB�E�<��T�$hy��£>���i��3���t�'*���gV2P�"�'�R�'>r[���B+\�7+6���V�U��}��F�J
k������I��Mk�\����'����?����n��@	���R�j�+pM��?����6�J�aw���wIe�t�7� N:�i�4�"D՟���%ɘ�[�ly�#	�5���P��iD.����&a6��OJ���O*�	�/0�
���J��D#d�6������^�[��<uZ�=����(�	�?�1dRcy*e�n�]�zV,䣴@�?iU�yKa�!Al���O��;��O�J�J����	��֝��M�d��n P�E����ɛ#�$=0"@�/Lv��	�N�F�*O@%�	�'^p����؟`�1a��{nȝ1g-���~u`C˟��Iߟ@�IPy���"�d0&�'G�'�,�����l�tf��7�� �'�r��O$Y�'��'�z5��'�PA��C*V��}H���WaܑR�n<�Γ5N�J����0;4l�-�q�t��?� ��q�X]�͙<����*To�����O���OƠ���;yO^������O`�ɼE~���e�w�p(�p�ǧ
^�ą�/�\ CTB�<)��i&j���d�L`I�J1<3���s�O_�̪4B@L�4HJA��O��yg�i*��;�~�͓<!~Q#r�aVn���a����d"W�N�P	t�_� ����ll ���	ҟ��	�?y�#��u��=;���8�����
�u),ܗ'��Ium�)c`2�'��O�\�j�O��N�_�
B?j��,��k^�6u���f�i�v�[��O��`�X��� �k߶��C��%���8�䑥-���"OwӦ��Aq�(��OF��D��@ERBG:		B@�Lۯ?��T���v���)/�(��E�'���'7��'��8N��eP�L2�L �Sl�R����)���䟜�ٴ�?	K�q~d�<���M�t�  `\���K${]`�y�J�4A�u p��_�~	`�Ɣ�<i#�C7!h�}�|�a@�|W7�qJQ&��?�6�c��/c��6쉄SdL�!�'6B�'!�4$W�C��OfB�̌xԂ�Ԯ��w{�dq�E�o2�'��C�v#����'���{�d��>i��dׁW� ��ūh9<�#2m�
t=��'�%���ք�?A�'M�v;[w��Y�U1O�����~�i�HF�x�B���Z� �'1��y�\��:���^Y����?q���?!�`�6`0v��̗�^^Ű��X��?A����ˠ+��4��O����O"�I�1n�ѩ�G�.U��`%A���r��<��S�`ڴBu�n9�~l��\��'?�Ic�E:��̓c�RdݢU;��Q#+��q�L�<�^wp ]I�'���#\�<�DN4q�ज़�%� :��"�kY��?����J�e���?Q���?����d�HxQ:�D�:�,L@O��.���`-�9S#<ʓX��' ��h�OFH�'u�@\U�uÂe��Y�~����ψR��ʟ�f�E�'N�7+���'�
��$��o��<8��'*#h����z��0i_XP�@B��-��)j*0k�W��?����?��'>�x�ɟ���
��e�V��ޢq���d~>4#�',2�'���mT$����'ٌ7�u��G
{>\�$JXoA.��1�O�����b���ĝ@�R��'U�d
X$���T�d�yB�^�zi$Y@�➰�|ȸP��ɟ\;բM�E+�ўM�f�IBg�zͺ�'�yze�-򬕘��B��k���;i��U�!��O�$�OZ)a��CN�"�b��:�
(�S@�O�	+R��� �Of�$�O|���O\�����)v(1�G�9X ��)��X]��8�'V����

�]�vA����	�)��dؤY(��A���G��!@sF�
>�x��gd�	�39`��)� 8��lK�&(�p!c �3/��@� �'�",ied@���'�,6m�O�q�E��8�� {��5�ЎЅ>�j ����&�аzQ#B6lL\��2?�F��C�ͺ$ۘ�y���Q������A��[�#@���N��L
����	/��˓bRkB@�N����'=��'*�$
ݘ�܁���?F��e假YdȔ�\�Is쀧c����������?у5�Yyra�$�����#6��=Z1#ѝA�b�(�f�{�` 2A�O�K�&��	Ju@�i[1�ӣ$�t�����53+Alx��H:��e������c!��6�|ʓ���]��Ia��0�`��+%��\���%��'��'#�P��2���Wyޅ��i�,�����+�P0[c��� �������MC����Q�'����?���Z�t�#�%�1K��gC"���t%T]�`��q�ѷGR>�I�]�b@�¾�NC#����Y�C`�U�b�b�QLK<`�ʌ��j@�YI�P	�kP���ßL��R��$?!�	���i�ccLW:�Ж�L�v�4`�I� ��H�m!�	�vy"Br���ğ��d&a�YP��>1�X�f�*�����'��A�o���?���":8��XwHl#�8O��C&lme!�ퟋ\���֜V`^XBf�O�ÅF^}y���O&Y�#בq�^�$�O����+ln��0\�O�>��A҅0�|���O�˓m]��hB��	��L���?!@�&=FB�A���;��h���&`i�'H�ꓝ?��J#H��X��(���?�qK�����pMV'O�fa��J>6��0A�͛i}Ã1O@�0M��b���Myr�L�GO�M���R�W"V�8ub�:��DҞ,�r�8VG�Oh�d�O
���O �]�Z�Z#��>t56p�@J�� ��'?À c���?)�i������dm}��k���%C˰%���@toT�$��%B����S �`O�*f���V2O���3!��uߴ����O�Li2�k�?�6-s�]�y�	/V�����"wN<�DV��$�	ן��S�:'���O��ikp�&A�p��@��!l���Y�HA[Ov�0��?����Z%����_禉λ
�`�J�F��MX��6\�<y��49�����~B%��xݨT�O�*]c"����ڤɖ m�Ta�'؜nr��� �}���I�F�|�Q�6O�+a�<	��'<ܔhl�*��O%Uޘ�EJ�B��`��ʈ$7)�'���'��I"!���������	ȟKg 6g�}�T�\�(Ȝ��c�ǟ�)�a6?	�]��"ߴ/��&��~(үN���� f�a2�K':��G ��<	L�)҆�j�4x�( )�:=�v<O��
'�ߵQ����B��r��X&-�+��}��ȟ��	�I�$q�E�՟`���<����	?���6�b���0�������<|��a�	ޟ��4�?ys�Q~��O:xh@5KE�� ͘��2pa2����P�	�<��4'p�T" �Nb��6n�M�u����l�7-�V�tbT�wҪسB���X����<Q5�'֙�&��#�b�'��OC̢���ou�h�qg+1�@��\g4剏\
�%��������Iޟ���Odė'S�@i���1�4)���j���a�>i��?��@�i?�t���W�`�'�8��9r5�bc��hD��G��k�Q��<�FJv� �P�5f���'�����.�H�7L}��d�E5(爅����*հ���Ob��O����<��)P��@ �>ʴ̰�
�"J��l�?p�Pe��pz���'XQ@�O���'y\7�AS���1.���k�J�`����0/Vi�$1��+=�$$ITw��iSΊ�/��N���!h.�P�;<_Z�lR(L(�ʳ-�_�8�#!�0�N����`�	�?���k�`����8B���9g0}�q��+ 2�
F� ��ßX���Z�{�^��'9r6-�O&���	?@'���Ӊ"^�f؈��<�<��|� 9� � ��5lZ�?��"��+v�]�yB	�%��gkIP-Դ*���	�>剔��ПPx�"�!��čޟ`�uS�N�� �	����I���Y��4YLx�tG^�?+����ݟ�'�j(j��Ђsu�'�O��	u�w�H�!�U�"nƨXr.��j��	����ܦ���4<dx`+�'����Bl�*��Q�	��ֽ��d�U��8K֏��.{�D�B��HD�+�č�<�Zw��\��]	Ȩ�O���>�5��Թ@S��� m�8g^Ҥ+�p�y��'�2�'Y��'L剂z��Sѣ�#bi�h����R�����t�1�'�^7��OH<*����*�O9n��тC�L.
���gƔ?J�6�ٴ]p&�X�oQ4j�btZC�G�<�%���5_�*IrY��ڟ��ˡ�\,ah� �Ä�.Q|�:ѹiƐ��9z\qd��O ���O��iNC
��'�E8��W�j�j�H��{���0��)9����̟����?�I� Rпi}�N�B���0!_�_�4�^�4A"�'�I��'KI���t�����fr�NC�[V�	aa-��ob�CL��,�Tu�tSڟЃ�ŉ�0��$+��˓Xk�ȕq��2��'�DCcៈ�4�wc��S!��!��'W�'v2Q�x�uI�L�4Е'G"E6�����Qrp��v0�㞜���{}��'�R%���~"g�5G�)����D�J(9�E=Op��G��<Q���*�����A���ɔO��Ћ�\,��ߴV�(+(",E�5	Q� >sM6��	�� �	8_V�B㍐s�����	�<Y�R�=a��0d�&TK��� ���X�����9�`i�'�B7��O� ���P�%;Ҥ|�7���v]��kX4G�-ˡ	®X,H�ɤ*��X����%�y�+B�2�;;���;���4��h�"�ŜM�v����T�_/B�hv�N�2T�Ց2�'�r�'X��!�d�g�A+p�86EX�b{hA�^��@"K�\x�����(���?��SJ�^y��!c�\�"DY����ҏH���?��2��=��E"����(�*�t��u+�$�4�[RiE;$.����+i��͓$A��SB�Otp�r�Py�E�O�H&늶��i:�˙L��Sb�-X+�}[���O�$�O����O��t����d�2�?1��äB���(@Mă +�y�E��?y��i	BN����$h}B�'�mA�;��$�"���p���c.&X#wC�^O�]��. �y¢�$r��0���ibrQ��tޡ�L�!)��������r,C��&V&�3��O���OP�I�NR����d2� ȼ��j�bm&<�Ƅ=u���Y��'��' �,�RF�$N���'K26��OdK�O�� 3K4jj,�S#G�.-@�%��~bÇȈ���nɪ�uG��D�3dT�	t�'N�K���> �f		���y�+CB�Ɂ�?yHD�Dۆ	����?��T��`h��������ӂPA^���?(O�-�v ׆n�����O������@�
�S��z)�;3��T��K�/�bʓ�����M���iAT-q�'A���u�\W��jO8�򼨀̚%C�z��s`^�7|�D�	�Ѧ���%��<�]w����'���jTZ��A�CP�&����өT��z�ɏ�?qb⎋O]���	9z>}R)�ݸ���kR�u4y96BD�x��m�	؟��4�?��l�R�	��M���92���Ҡ��K�ؐ��l��Aޛv&�8{^I���ּl��,Қ'b����A�o���I�'.r�q­J�l���rB��I��An���?��>-�����?�����"N�/��Ɇ�v�:�"v�O�c�&AJ�i�o?�lȴ��>F���'��O��	�t\��
�4�y��4y��D`�	�T�uڔG��!=�&{���S�Ov �@�ͧ��I����]�@^�m!PڨC�B0C�D�(�˓9\Re�;0�1����.O��ɠ_5�̳�D�ڟ�!6�T�{6ny�@ߤt�@�֟��쟔��{y�$p�9��'�2�' �q²FT=Uv�
S$-�:,8��'�2��O�]�'~06͔����� �r�B��Bez���c1�Ր�eW�P�L�c<O�ѩJC]�7����OΖ��'Ў��#->d���nC�PL�=P���h�O`(9W��b��xR	��ٰ�d� ������?QCN�?ue�m*���?��ih�P�������s \r`��: �ʿ/As�$_,~L�����O�����%��g�.8�+*x��4mu�7�!�>�S�@��: �yp������VΤ<�5�'�b�`���,���'gr�O�U��+6�Tu�Dă�7!�]�sF_?0��I*���UeGٟ����8��NvP��'��� T�Ӄ#ĸ��u Ӈ"E�Y�(�>!���?	��`?�����{�'O�r!B�Hc���DkS�|����I�7����%��<ٷ��� �.�Dݞ8vm�'���dN%S��b`�[��n�2$�#8�T���F?9'����O���O�d�<!e,�s?�D0��w��8�d��RvxI��5$�"-���E�f�'���OV<�'��'�����^jn�&E��@,��c�"����+F��>b�'/�I��o�ҺoںP]z�O���o���r�6WX�E��s\P�!�[��j4aWf�'����CeU3��	�)��e��y��?-�M���
J�.QX)���o���2����a�����c`�ߧT�K�'�H J�'�RM#%I3����O���c5��*L�s�j��SΖ�#��`;�GI�E���iW�M�P�3R<O�!� ��\C��\�HD�.�?!��?aG�߀p"�R@mX,8������˵�?�������`1;$�Oz�$�Ob���4[Djq�S�
2 ���5jL�R�X����O����iy��'ݛ�%Y�~Bɑ�5>�XR��2�2Y;�k_�:*�a0���X#b(�e�5& d��޴����'��.E� ��dM�G���kU,ep�^�xW�8�#�K���X�a�'��+s$�0=��-O7PAA�⑆(hV���V�NAR��
�?���(���'�rMx�O�d�'Lp7��R���K-���x��@<N��l�z�ʬ���V�x VՁuoh�����L�<^�i4��)�ԟ �2e7M6��x��.	�|] ��i����Z�d����%��O4���O��I�+̖�D��i��glQ�͌&U&j�3	�RP��֟����?-JӋ�Ey��fӸ��*z��I�F,C�2\�z �zK���I��YHĥ��<��R�#���.�:Xw8B=��Gج4��	a��OE6ͩe�׺8�n�$�����V�xy��\��s�*�����
��?AA�b�e#���25�@��'#��?����?�����D�C������Op��O�Q��>��X���~� 5�c�O�Y����:�O��m�$�M���U��y"�y��Q��i�*�)ib��B�/�<9��&F"�
%Y�GL���Oe<���h���tF�7FSJ!�LX�hD&�#�Ӻy
����O���MW1���$���O:�dl�$�d�J�_��Q2���14��q���O&<uNV;x||�-C���'^p�O���CQ�D����ټv]@bWc˿#4����&�9x���oګC��ʑ`Fʺk%,޺�y�j�ly����b��#�Q�.GR��G#)\~����IN�˓a���\D�b��'�B�'a��O1Tj��S* H<T�W�Z�6!$9�ST���D�
,���	П��	�?%��`v>	�� �N#��[B�(4��& z����O���O4ԣs�O�l�����i�M�b����8H����M���P.�M��b 0�y"(ʷ!�_fpջ(Ox5�����)@$D6z�Q�Cl�� �zu	S ͹Q���	П��I���Hy�nI4v^`P��?O�`	�����A���8��J�'
7��O��&���p�O��$�O�}y �3A�~��F��*V�XR5�Qo�� �)�p2.��u9OI�4�ݳ�u�4�!+����;e42�3%"O;G��*�k��Y�τ9U6X}�I� �	�?Q����u����+�FǙ~�|��h�$Q��=����ϟ��	�xCWK*3�����؟LBߴ�?a��B?��h�FQL �ǥ 'W�]Jp��?[g~�	�I�&s�¦�SJw��;;<��zq�'��d٦�Ϟ��0p≐,X����^;���͓xnVuQ)Oʹ�����	��������@K�mI� ֩�  �ŪI����Izy�!��E��'�B�'��� M�U�����o�KBꎌY]~���	����k}�'Q�珥�~2��1$e��'�\T
���,򡑤
�.VQ�,;���( 4�)oڂw]f Γ�u׀�y�Ȕ$^/�]r����;��
`�>v<z9���hU@i)�a��?Q��?���?A,O��@خPtF��b���oعj���v��E��O����M�	)v�X�p��	������o��᠓����'�� �V�Յ���Rϐ h�f牀G�\u
����+.G��	�&Ekf<�ħ�(0�^U)2-ś4��V'�O�	��l�����O��D��I끦2� n�qK��o;R��a��e�VĹ���??ԅ��S�l���?)8�h>u�I��M�w�f��"�>t��H
��P�^�܉��?Q��]?����_�'�ܤ;^w��M���Eo��q��4��u�/H��dJ�3xF4a�'tR�O��	w��%��������!�,������7�8dk�� ��	����}y�b,e�ARS�'���'dp9x� @��=�t�ڬP�T�F�'��e��O��'M��'�}y�'@�᪐�B v�޹�,�8�tkd@.E���A(��0'�H$�McU�ߢ�򩘾 A�d##z�k�FF�
�l��w�����`�͟��	ǟ����*�z�%?��������P��@�*(@��w�U���g�'��]�ҨLH��	�M���r���'Z�ԩ_�3������-u�H�/���$�$)}4���'�HղC��4�L�\�	�y��t84���m{�#�(���-�I�"]�R)�=:�D�,O���	YI��QA�̟(�I��S�p�x�&R�i�<�0a�*�t�# e�Kyr*��
J���V�'*B�'����T�.���6b+2��uǗC]����LA�\p�O�n��M{��o?��J�65�V�+V�T��T"����.N
����L��M[��yRB^�c2�͓WF@H�/O̝�I�t�a֊IP���[CI�Ӷ��'�<a!�	��<�I�T��Fyb�͍]]:H:�'�k�-M��xZt/^"Ȧȋ��'�d7m�O.�E�� íOn�l�M�R��d�hiCLZ�<�Q�XB��`���	<
��<��O�/� �}� IH�ŭ|�&4���.��|��j�5/����aɓ�!a ���'���'0����I��O'FPH��]V"�<��ٓL];r�',�S��޵c�Q���4�?�$��U?9rǝ0���G�h/��I��#r��:&�<��`��M�� ��䮻X���'�r�$ͭM�0�Hn�&-t})f�����c��D�-O���I]�����Nޟ������󗫟F��1��ATZ�T����gy� Zl$T��'��'M���2B3~܀�-��K^~�:6��W.�hBX�੭O��m1�M��ӝ�y2�B`����� ���	� ��M�D�P�Zy�g������$�Q�*��溳�D���,������$Y5j���@�}B����x����	Qd�١#��@�	�(��ן�'�@�dj�ii�Q���	z�p9�σ6y�����'�Hv�����7��*����OZ���D�>셚'Aƶ)~�R��O@�cglW�Af����E�7�D�T�މ�_�M{�j�����_�I;�� �[������M�'�l��f���b�"�'���O�����?�� -S�� Cp�0'�ƽ2��]�<��e���OV���OX�i\�%��	�O��n�鼛��X�eO|9Q�/ �4��Xq��	�5������LY�?�C6�ຫf�U�~��3r�=Qk���fK�z]،c�'�L�����<!DA��D�ܟ�S��Djd���I$��a��	�=�x�D�u� ���ğ@�	ԟД'Z��YEkS�KTr�'+��Z�C����wMMÕ�� #�`��yb�'8��?��"�f���������ec-3�M_$	���FF�toj���=��%ye�¦�ru L�<�_w���'A�	(� 
�L��@�/��\*�ޟyn���Ol�D�5H�rg�:���O��d|�JT��yR��"��/����r��Otp��+�.����OF0nZϟt7K|���	�?�ȕe��9�\��A�����
�Ӊ,�Ȍh��M3��-!Q^�#\w؆H¢��O��Qe�t����-�d5�J p�o�74ꎍCe���R�'!����4$e4|Ñ��O��D�O:��	�S��|�"�B�ct�J��̳~�$I���<���H��T�����?����z0+��|z��F��pb������
��̸�^�dS�4A�v!ڋ�~�!N�(�(	��'���- �[�V5+T��):�`#��P�	����4�ȵɛ'�\1� ��<��L��$�8���4����D4�$�7Ʉ�J�VT�p#�<�"�'���'-�]� c#NK�q`z��>l1����ְ�
�ݳF=�p���M;��^$�'���?yܴ=ԉ) �5=��@{V�9�֍3�F/ BQ�G�Wi�>�ϓaĵ +t�7��5-��'i=�nݫy��fN=`0{��n0H왆g�Vy��'y��OalI"S����'x�ـ&G�dW:�/���A��#��'^�J�%T��|��'b�r�T��9���A�u��횗�&Z��q���Q7t�)�'7|�8d�:����O%�=���q�0�k��
�g]"'�-sٟb`�K1�W�M�y�8OX��t�<�A�'n�I�t�Ԍ	���'^���b�+���,ڄ��doZ�4��'�ɯLr��a��{y2�'�����:�&�3`��otԬQ�K�
z�4��\�H+O0�$b�*����O
��E����d/��cy��3s��-F����ɬb憨`<�M��÷�y��*`8�1O�I!�&�<Q���s����c�ăT��~�"cӍPz���'�2�'��'$剺N븜�Dc�p�` � �V0ɲ�	���U��ɟx��4�?1��Uj~�#�>1��Z�*i����;O����Ȇ�����}�>,@���;�y���<�d˂C��}��R�h�?�+p�%{B\Q�jI�ZT�y{W(o�����D��(�䉜��X��埄���*QV��O���,�J�x���CI9�P��kA�~	���?a��귢�������ͻ,]6#4`<*d>�*�ÓhM��I؟ȫ�h��X�ai�
�4����2�Q�s�YZ%n_�`3�A�ЋĔl�9��j�,\[�
�����q����j�Py2�O�٩@�ӓ"���� �:��XHS���;6�x����<$R"���O��d�Oh�\|����Ǚ�?����?��i�.eKy@��aDZ���K��n��\�I��	ԟ��I�"�@��2S�
!��c̻n���	�	���%����$h�䔕"�`��Ul����t���;3����qډ�@��[�J�8��[�Z��R��W%=��'�b��$0� ���D�':�0O�m��셊j��H: �wƎ���'�ʐ��g�wvR�'ʨ7m�OR<k ����Ӡ;���#"
��QC^= D��.%�x|#D�ǿ[Lƨ�I�@�u���Ժ%����y� ��A��P���� �a�<4<����ڎ(��-��mb�bR"eG�=ڤ����'��'�����%Sf� ����&�\Xw#D�\�Q�La�m��`�����ǟ����?��]yb��+Β�ұL��EQ6�ʀ�Y�1pN�UH�#sӮ4�-n���F�I�#0�ө�,�@읁��ձq�S�G���]	���q���`թ�B���jT��*�����d�1�5)Gm1�a�L���'�T9 <��'*��'�P��I1�5I�J�	En(2���,C�H�Iw��ECƐ�	(�M��
����'���?a�#(�1�,����EEAu�d�%�qn= d�=P0͓̄= �h0�}�7���Ђ˧r�󎏑]WhQK�%� z�py!R&Z�����`�p�b�'���'M��$�5�ObEB J��$�2�;oae�M�Y��'��4f�`3P��`�4�?��K?q��
O���ZV�ŜS$�؈�$�=WqD��F���r���M��'(���Yw^�	!�:O��ID�˗B�X��f"F�f �M8��7T�*q�`�`�j&R�X���q7(�A�R�?q��?飬_�o!�1���k�Pԙ�l�?	���DϠw�8���i�<9�����bD�`�	�(�ց�$��pl�+O@d�'��6M����	�jP�<�V���_���ӄ�>`�'͉6�R�%&�V�\�a[�X��'l9�de�!����O��� ��^yro�(fԢ�2c�&a�L	�5eY��6qY>�{E�Op���OZ�d�O4�f�6M�c!/,av�`��r
}���جk	 ����?a��i�(H��D�\y�'�����V�#"�}`kYa@��i����^(%�=ch��y�!�Φ��_�Mխ����l�.^g������9��4�C��9�M+��'vt�7Ǖ�c=B�'�2�O8ƌ���?��f!i�\ sgJ8]�����$��\kL�O��$�O��)���\�;��V?���[&�\�B�n��p���"�R&|�d�o$�����C��LhP�?�{�!	ݺ����R��KG%2^��1��4^�� A�'Qp��4D��<�bE ���џ�kc�ݱ8Z�8��D>F1c���.�8`��P�jZč���d��ğT�'�5Q'� x�ʟ<r��B��Y�I?_#~������tS�/1?Y`S�tY�4v���;�~b���
�ʔ��@�5�jT�0���B0x�ٴ�y�ι
�0�b�i�vŠcU>�S q����H��I���醮�6q���1�&x�����?Y��'��Q�צ�䧴?1���yҠ�?^��D9V�|i��{tK&�?�D|�,\�/OxlZ���jt�!?���z�J�x҄�7:�Dq��C�R�-Cè�LJ!��v=sG�&�uwE���ݺix-0_�MSs(F(5
�u�E�*��!���O?_i,�3*OT��	�
v�y��ğ��	�|�ӓ" I`�h�8
p�,���	ky�l�7�x��[�p�	�?�S �3�A�/Kb��dO�#i7T��e�̉ ��IğH������	/!��`�?�!R���|��M2W�%?�e͜���l��8v�̓-�*e(d�z���C-�Myb��O
a���;F��	���ք�1�J>l���O��d�O��d�O@�����K���?�͖&u���3r�Q�u�B}��M0�?��iJBb�����l}B�'���=��!�i���p=x'ڳb�Y�MG/t�=�uI��y�ӊ%����e Ӡ�X�D�a�J����K�4��F+�$���2����h�h��?����B*���'�?�#��(ò����"��e���R��?9��?A�VI��.Od�lZПh#d,���jBLG#,j��f�˙]R] 2��+����k���'�����%���g�0��.<�����K��})���7���FC(K��ꈗI�pʓb���M_L�b�'�b�'r2<�F�opl�C�Wr��#t�'�BS��4h<1���͟��	�?ɰ���zp�0Z�iW�H�)��
��qG����hجOl�D�O
)C��O��!��*D�rM�?������JB��Ge�|�s	 `R�L���l��W�N�J���Wy��Q>��-3NK���q��k �B�	4�^q)��ϮY�
\���� b�t�>I��������69�L�V+�>�p�(�L��?t�eb��7���_��ܨ���Y#��cႏ (ؕ�I��,r�#B�-,e�HiAP�4�,8��@�L�ۃD׈D��xb�b��@;\Q�%N�6BZ@�,�>J����Y�xhՍA��hr�"��E3He����!G~���蝼-�\����F#T�r0eE?w��{H׋Ig�Ar��79/��T�*���a��L�9m�|c
��MڞyCtGP=z�4�;�*lf�\ٖ��/M���V(O�r��%�'�ȐcUt���LL�f�"h!��n���毕M㜴�6��|��IA���W���qwIG�R���`4�	R�F!�e��y�L"��� \.�����,<�t#@I�t�@�b�Û�"Hyh�"�$4�h8�TI
1lOPA8��[�U>X�AL��M�f" �fY��Y�f�]� �"%G���yr��<��B�	�,��S���qEX�����t�Si���$�O��\6ͽ<	�LJ�o��O�HY�paJ�~��k���0U\`���'�.��~���$���?���[Ӯ�Z�l�TA܎'d��I�t��Fy�cY=T��r��꟤�;�k�:>�>a���N	c���(�ڙ?�d�Hw�)FxrN�=U�r,S����� �?i)Ov��4Næ��OJ�O��W��ywl��%���R$�2P�(��@������d�y@vQz�R27\�����q�`�4d{,7m�O��O��iVey��<�?A#eWi�)CqIS�v򉳃 ���yRHLF� ��9��!��,J�A
zP�i�*0�b� Ҥ��O��D��%_fi�'���?�4��*)�ji!�'I#NܭHF��K-x$
ߓ�?	���?)��6��z4�@�G�b�yħ���?A��p��E:�[�D����O�����'6�<��0�M�3K��8���8{��,O��@��O���O�ʓy�H����
}#�<�⌘�g��j���i,�I������O����?1�'#2�ab�B�8V0�Q�N!騬+�B��T�'p��:�H� ��n.�rF���k�6��$�2��ΓO`���ϟP�Q�Rn�d���g�? B�UR6"@L1	��Ծr��p�Z���	ǟ��Ijy��݂1�N�����-K,؀ɤ�A��������O:��I d��D��x��)�'Zp�+�o9�r��'�nB�%���?����d�	"�Z�'>}���?�A'���0�m�Fk��0���C�eh��n���S���DQ-{�)�ԥ�":)9��lQ����j@�M�(���$�zՖ'��m����&����D�QF����"C������p=Q���AR�ޱ�z�I��������"��M����?����T���&�t�ġR��4Y8�Y�!艈��Y�L�˟�`�j �h^��<���{��%[���r��@ �F�t3G�i��'t"�#3..�H�Γ�?i�e���@��4X�&ѳ�n_?,���C�45��'fB�'� B�V�%�N�k��@z ���'�` �G�>A ��<�-5�y�Ӽ��A�ZV�=4,��@,�Q`$��syB9\O�V���Iǟ���Zy�ݦ1�L���)�!��k�ǖ#~]���>!����<���94ܨ��?��I�,�A�e� D!F+*��q�.Ρ�`%�T�	��	Ky2,No|�)ڞ?�����L;I��XaS��Of���yR�'�����j��?1v���?	"n�x:!��M�p�JƎ���O �d�O��2��X�Q?��	�b���#nN�W�0xw�ߧ;�0m��̟؈���\��G�Od���$�b�\�E�R�B͆M� &�%_\(֡�O���O�˓E6|��Y?���˟���-x�4��EbDS"���wlI�\��������iע�O �DY��̻(zj�"%Y	�t�3�U�g%F�	kyR�_`.�7M�OP��O����s}Ҫ��I��iPW�۶j�ZB䍞)h��L6�'dR^�\��O���~�i]&F �d�Q����ɡ���L����Mc��?�����gY���#�b��2����D�P�"�*(��T���M���{��Bd��L��)�|*��S.Х���bd2��$��t���:Ѳi��'�R�K&?�\�b�X���?af�	g�<[ï֖2�<��SG1�:L����NR)�N~:���?�5��$�TlsSIi��X�Ya���?AJ�I�I:#�d�I(�����]b�� �'a�;ad��R�Pײ�]rfyL>���?������Ԭu�s��R�d��Z��PmMy`�yy��D��?I��B^��|�0���Ϭ
PX#�Y2!�ƴ����?	.O����O���<au�Q�.3�tHЌh,Mi�,�����L�y·'�?q�/zL`M~r*� �D�O\@�rq��9���K���2S�6˓�?����?�,O�t�"�y�S(&�~|`�%xF�h&Z N�n���ן��滟l�ƾ<ͧ�?Q�Sj�B\x��T"ځ<���������Iݟ�'E&@��o>�)�O:��(r ��Ѹ�{�F�p���#!hZ���Q�d��	�?��	����<	矴T4�lɛK>x0�	�?A-OB�7�Ӧ��O@B�O@��|���M���|c��' $,��{y�M\%4�r��9O�Ia�,J��L�=h��R���{�r����OR֭B�I�	�p���?�S-O����Of�)9�n 4Z;�| �������'�p(S�'�R�|ʟ�I�<�����S�9o8�7fS h~h�	�������t����vy��5���9O*���*��H�KK ��k���<v�[��d8�Ɵ��W NT!UC��,^��B��]�-hLU�I֟t�a�Rny�����1O`�����)<C�%��K��%��|������Z8��'y��'�RQ�@�7KY4X�����զ���ˇ̘N�|�-ObIIW�'*�#ۑ��y�cF6��TD�ԡo\ę�����'��'1r_�t�I� ��̧%5D�h���=a�>�Zè�)g�\�I.����<A�@�����O��'T��u�*#(Ϊ��f�=��2`�ք��$�O����O�ʓ2������$�˨2X��AØz���̔�|Y"�'7���'��\�*O�)�O��ԟ���C�#D��K��R�s�'BP� �	�Y���O��'��Ž}��p�K���3�F�! �e �'�W�O@�����I���8����@�?�8iѣjy"�'S�iq��'���'�B�O�i��M!j_AÐ�U����
�35���I�<��O�3_�#<����(�*�>oEL-h@�<���f�'ȼ7F\�A�	���I�?)0-O>���O��y�BcNJ�xԫ���3�"]��'6$�p7�'���'��Ic��'��)OgN�B�8����ي.o�6-�O@���O�q��P]y"H��|b�B��D��m5�@�&\4�a!����v���O��O*��<i��?��@����Q.��� ��Tt<��?���3<B�� n7��O�4�Ә?� �@R7%���"e�:�D8�KB�	۟�$����Iy��'1`�S̆3�x�R�:u��MI�ܽJ��I1	d�\�	�<��ε����OB�	�A",GAX^��h�㏘M�x����1O���<���O����O��Hz�?D`�sGj�M�P*��j�@����y�fK?�柸�Oڪ�jSM�~d�9�[+(��� ��	?%�ݟ��	����'8�Cp&�~b�V�$Bu�Z>��`�#,ʰIK�9����?) ���<�4�V��?A�Q<���D̓5_�y��i�T��M���ƙg�����l��Ty"��/)6lꧬ?1���rFd��u)�9X�/׋S��}�� ,qդ����A1���?�(�|~BZ���{�? �-'\ L��2E�")C<��b�'p�ɴVE:���4�?����?A��%��	��5j̫�68YG�o����'���6�ǌ�
��D�O�˓&P����V@�
:B<�!�hǝTQ��ra�'�Bd�ԩsӜ�$�O����x�'Q�5؜'=`쪔��9b�=��+�{�(��'ȹ��O����u�|B�On��x$h�8��ERD��7���Ҷi���'�B�a���8qV<͓�?�%h�6gM��Ӫ�>@�Р
��5��S��?,O�ڇO5�	�O��d�O���p��zr���p'ЍIs�!0#��O����:���'}�$�'����0�y�wz�8��q�ЭJD)b��	 ���?ҍF�<a��?����?I�����Q�g8UX�!W ����ԄCf@B䃌E}�$�<�y"�'w\;�'L���'SrK�!�2��
۹/�h"c�\��N���'���'��'�2Z�ty�����d�Nq�IR���(i)�aC0�� C�h��ɲY{��I�?M���`�b� 4��Z0�Q+6@4К�JYny"�'�2�'���D ����f��I�U�а�ƒh{z��C�Y�-�X�D�O
��Q9O�eۥ��O��䕘W�i>�Y�*))�M��B	�	��SI�0�I��'aJ	��$�~r��?y�'Z[�d��^�3kZ����Ƴ(�,40Th�<1�(I"�?���Q�V��'��I�+�n��ȊR�ٺm[�@ 3�ȟ�'v�J�l���D�Of�$��P��'�d�:FiS�!���`1#O)18��SL=R��'_,�`����1� �VA�AƄ#"�xId�d� �ɂ0&&@9ڴ�?9���?Q�'TD�	H���ɚ��Q2j�(<��%	J�%���I�c����DΆu�1�����
4�=��쎂22�!�F56�B�l����	џ�H��_����7C��D�O�|��D�a��0HT�\�d�Ux�D�O�˓��0�I~����?9�O� �kR�o8�\��Դn��:��?�bNT���l"�Ο\8�m��̻	� 2v��4�Ht�)��'ʹ��'c�I���Iן��'����M$��P`hț=W>�b��د���G�����?�����<y�'�?��A'8��IG�<��4���b�fUc%���<���?���?�������>���ӹ�=�d�3c�p"rg��'i<���+��$�O0 �;O�I�O��$U"|�d�fX�6n%|_���ga�.6;0���O����OH�$�<�Q�T-�S��o�=$� ���%��N�ןX�ɽ�2�ɼd��x��埴XA�<?�'6�X�T Ix���$KyQ,#��?a����Ć���O�2�'>��ɾ)5
 AD�)j�H�!A�&L|z�'A�8Pc�'E��S�OJ�0�h�p��In��YwC�J�|���<Qԋ�c��6�'���'>����>�E�R� �@�`HK�.�I2��z8�����?��j��<�O>�B��j�i�/]4V!H���7��zd�N���n	�daj6��O����O��)�My��5�?��<:�\y�*X�JT��Y� ̀�?)��o�'y3�yb�'#����j�(:��P(%��T`�in��$�O���3Z����'��%��?��K.CM��J�ᆦ�-J�i�&9��)�����  J~b���?a��¡�Ɏ�� )X��C�	�jMi��?�񎞘y-�	;[�����O�I�R�?i�'��<m�ƽ@5��6�4$����[y���y�P���I۟|�ICyB�8[�:�1RG�+@�H��	F9L���ǣ<av#e�`�	�$\�'�?���z�j#�X�C��%BǪ�:l|�u:��@g̓�?����?1,O�[S��?M��� ��ޜ��dU�;������a�p��@�O��DN+,�ʧ�?Y��j�TEa����8���ϒ�*a��Ě6U*�-O(��Or�D�<��'_*r��O��m!�̢6������;:� ���'3���~��@�?���a"l�K����$��H��r�]�41>C�!� sb�' S��S�#���ħ�?��'{`�e�v��B�L4S ��@�)���Gm?ɠ,�p�I�oD�I`�I׼[��ʽ刼 ,ަ	�����ןؗ'~�͸�m|ӄʧ�?��'��$h���v�N`�
Z&���C!�O��� <����� 9}Rpl2 ����lT���ݪ�?�E���F��V�'��'��T�<�ŋ�ڟ��cO��AP�aH�IB9r�e�W�̟�i�hUƟ�%��Z7�7�͟�;��)0�40����Y!���p�F5�M���?���!׮ jqZ���BH�OD���~[�DI�B�f�
�'�2��g�O��Ox�	�b'���O8���O��r�b��dBJa���V�K`Cd*�O~�$���(�'~����?���H�][��2rƌ0M���c�\;"k��9)O��A�;O���?���?*O�c�����Tɕ4W2���썂V�`��'>����?	a��<y�'�?y��@v�x��mR�
a�йt	[
��Pm�����?���?�(O���!��?���n��^%�&m��S���#�a{�d�5O4�Z=���'�?���'� m͓b|N���IO�"٤�PL՜-��-�+O��$�O����<i�h�)ƉO�"�K���/yb���5 �4jCrt�W�'I2'T+�~��,�?A�5������Q�X�`��$,��1B$���nG��'p�^�4���Y���'�?��wK����(��@cb$�1i_L(j�(�O?ٖJq����?��Ik�I��ب&O�.��),a�h0���̀]T�m�m���'s��!�<�"$ޜq�|Eqےw���q�&.ݨ�	�<Ab�ӟ��?��^8�Ep���h@M�`���)F�'�H��'4�'���O�R3��-k�O_@ȩ�?J����A��QĠd�";O��(R+Ą�O1��d)� i��".��\v���j�����p�Z�d�O���%'��'�����?��J�V<nP[AӘ5�&�:G�^1(�3�R��֘'��'����6p�@����u���Φcx��Iǟ��pD^���$��A��'v
aɟ2� �+�2{[RdB�o�+]kʙ����<	fMr��/��!ZvH/6��ݸǅ�Yq�Y��
�H�J=xa,˻f�HPH��D��1��Wڈēv�'�Cu�'�]�����Jf0X�D9"54�+Q-�/`5D��	Ο��$�D~���Γ�?���8ڬ�����K��G/�?�fA9�bJ���y��'��|"ͅ�2��HR�ώ#�2\yǩM�LR�T����O��ϟ���s�S�v�$;�^�s����to�Z�kТ\��|��q�v��y����'@K�-pp�N[>���aِB���'����1�9��/r�^uc�O���HY��n��G*Z0	��iv��p���1hT�r����qb�x�u�%ڗ{�"u�S�E�6��dkG�]�Nz����\���LD�Lp ��#"ՉG��աЯH���ŅV��Lɇ&�Rcv�atK�T߼|I��ʑv��%��`��T��e���ĉ)�V�4��edF��D�'�b�i�yH`N�!~QJ����c%���3�> ��a��i�y3�O�d�ݧ���3O?7�ĥ]Hs�J�k�"ِ��·4z�v�N=?��1��+|��S��MC��)8����� �6Kv��H���ڦ�8um�Ot��(?%?�%�h;Uk/"�u��ϔU7jq�"O�y[���"LZ��d!�b8Lͱ�|b�e�0J�$��?��	�MO.e�7��S�tL���>e�40����?�C�F������?����?�f��e[ܴ�M��aΰf@�h�
H;Y<��'#X�Jq��a&���g OԌ����50������И{�<aK�Y��hvاI�D7-י�0<IV�Һ4\��r��C�]�w�}�F -�?����hO��x�Ġ)q�Z0-�͢�/3D6����!�?�������,۩G�p���NH�n@����Ov�<Y�I_8H^�Y5m��@��`0"��\�h֦��?����?��sU�Q���>�?	�O��	�$b�F��#�S>g��� �LM�:����ӛ\������x��{�G7p��`e.P?!fN�[�l�	rAl)j�g�V؞p!���O�6�6~wν�P�Q�y¢a@|nN�G{����[����G�I�F,��ώ><C��?����E@h|�p ߧz�]z�鍇%�b�I9|Z�eyb�<P�����?����<�쓪$=Б��k��1S�A���I�H�j���ݟx�	�vpL��D�JU��]��I_*n�T�E�P<JaI��=,':(���D�t����_�8�l �|T��:P5��	��Ӂ'�Ԁҕ�C�'������?��T�
]�IYc����g.M�����'�amF�S��pw�|Ju�+����[������Y(��RP^��c�
Qp�(�
�)E��	�𖀂��{����y����62�'ě�&��X�1(Ң�"��(0�J�${h"��6'��M���O�ԧBë^'��L����M0:>ܔC��&0�m9�+��M��A�E&ր�Ԫ&�)���)��>S�~�s�_BvRp8D�y�Pp��'Qb����O"�x1�xy�"COlYs��$�y� \�p~>��-�uw�iB��W���<��$�-R�����O��1"a�;Dq��BN�Y�T$30Eȟ��	9��hk�����P�	*���Nڦ��`���P�����2Z���� �>ywlBdX�<x��ߡq��F��3��M��f�>��j�iX���Cʑ�7�I�$<=������>�D�܅�	~�x�$M��u�����$@�L����ǟȩ!���]?
u2�)��i6Z�a�ςe���Ex�'�hO���C	Ӽaꐅ�u��0�D"O��سJB!Nܠ��a]ʍۀ�'�(8��)l_L�;w#҂:f�}�*�B1��5�
���]�LE20KLX�$L�ȓPF�%�я�.
ݙR��7=xy���dHy�t?^!�� Ʉ0���i�I����rfh�1WU$��ԄȓB@��������)�d[�0]đ��U�H]�%E,~	�3�E�<�
�ȓ1s��ѳ�C;8	�����^��i�.p��%qB41Ӫ3	W�t��++�eb��ȪB��[�J���M� �A	V�F��ҁ�%��1�ȓpP��r$邨�& �(�''Y�ȓ+�Ti�׉��q��(�L� ?���1��`Wo�Xh��a
��Ȅ�px�Q�D"T�OD������%�p���S�? ���]f�|����t-��"Oxl(��_Qd�щ�L� �0"O2��po�q�nx��K��Q (�"Od͛���V0bQ�!�� �Z�+""O�@RK�= Ҙ����IL�A "Ox��i�
(~��Ñ$>^��q"O��%�:��TX��D"FFx)�"O��3uC QD�"���C;| �"O��t�F=A�Bah.�2X%`�*"O�M�v���Zo�M��,^9��"O�����m�Ԝ����4V�1�f"OhU9�N�:dA!�
L/~Dqa"O>I؁��s�z�1��8$XL9�&"O�š���YT�xF�FP�"OFm���Z��	�w@]�RK��Ж"OBD�	��ebzeC�T�!�!w"O<��*�Uf5*��4d�c�<a@ �t
x�C	��)8Rm��B�`�<	�M�E� �\���h�m�Z�<ɤ��� q8�I7@+��5�%�U�<r#Rr���"6-^#�L����S�<Y�F�N�Ĩa��;K���P�Ir�<�D�ɫN&x(֪	�yb\|��aYBy��X*'��OQ>�ځ(�32BPY@���j<I�2D�$2���a@��q��3+�4��1�3��4dQ$}x�4��ht�Ӌr5"�p6�=7�6��	A~�Á(K��\h%&Z=~M����;���dT)UЌ��."�n0�mS#2���X�2��/u�Lk ���Dµ�E,���}a"O�
 Q-i��r��һZ�b9��]�D3�e�f�qO�>5��m˿,�Fpa'҉y"`���"D��Jq��Fz��$�K�m�0o!��	�?��)�ϓv�P������.`z�P�D����?w�V��{�H�Yp�.~����l�<1W���p׶i�b ��}&J�)��F�<�gG�r�2q����3�>��SF�<�s"	,9�}*�lZ"W�dP�#��<Y��x����NM�d&�³��z�<����)�5�$BE�=M�PzC�p�<��hׅo���ǂ�	"�h���mh<�����S���%�:{��� )SI�+�'*�ٴ�
eBd(WeE��D�`�Ę� �*�$�f�jq��Ѿ�b��u%T�4�!�D�
;���:�cP�``Z���?JÉ'	(��IQ�S�'-n����މcH<�Av�� ^�C��;1���9ƫ�na��@C��[%��=�.����'����+��9��+B��4����'�P�-�;,)*�xun�f���J�\��I/\�&AB�1Ύ��'��l�����N?`1�		N>A�\�=���������Qt�<���)Ƙ���>�)�S��v�?�!�?�}��FU�M�2dYBiД�"�z�HTr�<A4	]��M3$���3���i�2C�	qe�	91��JұZ�%!X�B�Imu\���C�%����q���C�I��f��力h���G��&Q�5`A�d
t����ּ$©�gA_'2C�0�Gb��T�!�D�94�M��K�3!��d�Aʧt�tز3�5j��6Dڙm >L�=�~�#O,Z�5
��(�H��� �Z�����G�Qf�	�.WT�@��8o7Ј��$��x�J>�5$V�&��>�OH�A�&434���撟$ނA��D��j�6ʊ����0I���R�jͭ%���%,[�C����@�5r��b�
 [��~r��s��|��ًLކ��u��O�j!�{"hB$A:���%S�JD�v�v�E��w�vI�ւ
��V���!�+_����� �,�$��n��(�F!*�YK��mӖ6�۾8D���K�F�V$r� G[m���|�R�m���_.a��;'�Γ-/����� }�"ܥO���v+E
��6�k(�h�&M�o�Vd���i�lE�&�I�i����5bUt��Oʎa`�%C)���DC/�x�PZ0)�\}�w�! �,,PW*�(����uLԴ|�	�� ˎ����R���3��(aBPFx��	O�-it![. ���U�O��F=�$���2I1)�vS�'�6T�f��	�u�H� ����$���́OCv�p'��nn��!댳z���$d7�'!�H��Jِ�8�*$D��X����kK&��q	�'����ˑ�2�*�����/GE����~�|)��߇\���H�2���s�W�j�i�E]���w*��W+_i�"\�"]23Py�������Px!GU>��T��lU8~�h0�4	B=� !(�5:�^���̇�J�(ܧO�>�H�Jۃgd=rs��!9��ٰ�>ʓ;���5p����E2�x��Ȣ�p�)AC<?��D>����{{����O*t��C.ْ2�$�#�̠���jgMM��%!K��|
d���R�!��S	7Ԁi�3{Z17n� =|8C�	�l��-'��ea���5	��I&|vp�"bl�t�Ʉ&��C�֐a���?���D�7����Y�j�2�x��w�@MZUI�4��c�d&RH�a���E{|*a���i�8��gAgy��	�{��C'Ә]|<��K�-�#<��@42� p��.�'�&���K)���y*Ě�&��Op5i�Ȕ	6?>E�Sr��k6d	7U\��	4�ݛ\Ѿ�"u��`O�Xk�+}���K)Qw��+���8,
�9[�d|5���fʏ�0�.B�	6n��9"�^�I<e��<�X�	#P����t�ҷ2��	<G������$^)ֶA�X�c�*��@p����$�4�3��	j�6U	AL�X��1Abǔ� ��i��&��~2Ή:�*�g�|�O���'o&xg�·�Zk���q=��Y���j,l1G�6�RcH|�2��!{]��r���VdS��Q�z��O����	��6��$%2&��6%G�V��Y"c	�V�BТ�j�0Hah$�S��k���Ic ��Ln>L�I�ŐK:n�V�\J�����IIF�h�(<�� c���W����O��1F
�'-�>�;"B8�R4F	�dv�ӧu�X$j�v(�q��?5��Q0�̏��?!P�D�N�$M�G��Np��b�"�:&�S�zq����f�&��n2}��I`*�� ��=���S��	.Uޑ�{!�مNI��P՞��"��&�t	�AJ�i�Y�L�%���a�o��<�6h�k�y`B.�����_�ArP@B#lm�'���R���i�'��5�Ѥ 0��F�~tؓ��6::���勊#�~�2&P�:r�E���<������pk�Y��[���b�|�1�O.�T�Ζ����RS@ҳ~�‫r�dy��,.4�g�|4���J�M�!����?	v�N����� ډ4KZ �W# i>M&Q���@��0z��a�e���P?廡k����� �tՁ�e#	D�8�L�0΢?�u�Q�,�O��B/)�8�h�)q.�d<^DN8�rkC�I҉Z!��ZD,����S~����a���լV�:Y�Ũ��~3�	�sw��q�_�<L�R���j�'
<s�!��Oƽ �ƕ�r(ҐKUkeƅҺMK�Ù-����j��c$��":�`��4>��I�G64
 �
�0}�� ?k �I�B�(�ڌ�y��P��9��FM$�r�AFg���xB��S����')[*6�:�#pBC�RIx�����?~���r�ø !8�b5�F?����wi*6��#��V~��}a�A�{f1)d�|axbn�:	@P�sP�!S����+I=z���!���F+��Ka�:O�8 �H4��*�"�9�{�!X^�FB��μ�33���ā �I�ǆJ1�:+1�©E�P<@ @X{n��#_�?3��߻���9k�BW�����O�7M7�O�\��e��} �e-�(��0w#�$iZt;��[�N�r,�p5�F-��|J��ڪS ����g�q�V���Xy�U±/�z'�HR).�x�&㚔�{b(W�KU�T�D�({sHQ�n|� �*W)�	ˀ�z���/!̭3��P.r��,H�W�����؝��
��
Fr��v�^7B����D�W��}`�O�r��Ռ̈́�^)��J�^x��k ���/�"� 1�ԱW��G����n!d�2��I�xj����˖w�B�Х0tz�-�9��J Ic��7/�?CQ\�B��U�� �D��/�u���G?v�P�k��yE�D+Tؔ`ʘ�s�4��~�%U�EL��і҅[�u"Sm_P�$Lo�,A�!�X%5��Ɇ����چ(r>}Nћ�yg�ܯ#��8[�$'/@�-	D�����x�ȅbU`]s&׫A�l0�O�t/u 喴6bp�"1���q��$
wbQ�cWdY�禑�H>�ׁJ�ii���0̟B���B���/O�,��!�*E���b,@�<?�}ѳ�D�`|aT��	/����y�'��R��ȓ`vJi���#�d%��y��Z̟ �1��*tΈ,!6ԗ-ݤ� �R� �9$gǆ'pn(*a��7K�=)1"OP<�6	' yӲEF � �1�3m��d�QA�,Xl ��ҞB#R8�}�	����[R��镨��E�\IV�F��xr��/-��C�:=�bL����65j.�r��ڿ6ǂ��C�F$hۚaK����d����������\���(�M(<O��	�^��xMɷZ\̩ط˔)P����B݂=�<!�d�
}�N�
���့��8+�D���Դ^��Dx�kP����q�١qW�1�}BH- ��b1L��gfl�:��@�<afY�bf�T�t�P�C\���@=Wd��H�fϗMr
!0�U�"~�400�Q��LȜ&N8|�j��q�d&f�xSR��Ra�j�a�`gX�����)+"����Ut����=]�@ bsA�5B�a|"���(�9�n*:�L�:Տ;�2d���/S��S�'d�A����3���hB��:A�I������K0�X��/��(��d
��*	<v�Hu-�FoP�i"O�$��/ѭȅcQ&V�mR�ݑRj��ɒ��x�)������F4]�H���O3�(�D(2D�bȄ&V���F=u%j͋�ð>@Nם&2�#AK><O��pԯ��sj�+�M�{���9�
OP<�B��8��E��gf�	��[�y��-)��=h���Sh �;S���0<Q��!���j�.[��Ez�
�!q܆�~y��`B�s�h�;�EG;\���'��Fy��)�� �rT�C�(���@C��;7�!�d�]'�`	9rx�ݸD�y?�'����I��|�S��ڵ_�|3VN�=܀C�I�>I�EBsO�f�����	z�C�Ɉ���Sd�6��E)r�N�Q�RC䉭z�ᖡ� u;Qg�%�VC�I�LHU��F]7J����@�4C䉏sİ�8�왏����ٟV�B䉈k��p+_�x��
%�Bh��-D��h�%,T�Kre[�g?D�(��X\ P�����#qF�h�T�:D�s����y@��B��. y�I'D�����T>[�X`g��,,�0��%D���$��+(j����Pek�k@�#D��q��~�1��a~�dz&�>D�|!��E<�I��I
�r��6n1D��5�U�Ġh�jc'B0�pI(D��sã��"���C�+	,< �P�4D�$�Eo�cZ��҉��� s!�6D��CA�R-Hz���r�I(��8Y�h4D���A�Y�\���ć���I�f?D���m�3��-��f�+ޡQE�?D��/
H�8	!d�*�� 4�&D�L1�I.W���xb�Ϥw�~�!@�$D�̘���[��6 �&H�(�Sr�%D����U#<�[fK	..S�Ѵ  D�8X0�9�x`B`B�@�f����!D����\/`ѶKp��D6�����=D�,���H��RԉO�]���8u�)D�h�N���챒�J}��t��$�O�8ZQI��"Ke�af�v��l�7�]�2U�%��'�����>�j�#���2'̔��'Ҥ���Gc9¥���֘)�� ��'y��!!��d�x��aҭs5P�	�'s�y�g���"T�\����n������0�+�+!ƙ!��,k$�8�ȓDI��㓁ͲL��)'��Q����3k�$뷮A=8����W5sP,�ȓ'm� [�f��|7�d(f�#$���?Ģ|�vB[2��C�˲fXJ��ȓ^1��z!c��s��,kw���j����S�? 89��F������T]v"O��sׅѳ�\��7��/4��"O�%SǴ3t��@��ȡu_&h
�"O(d;�ըK��ab��L&��9c"O��p��Ҧ��L�E��9F%�iK�"Ot�pA��&TH�E¾@䨉"O�32����(0�F�V��}Z�"O��!S  ����a#0z����"O"|���	rL �K�X�h|Ht"O�qk��U�V�����V_�(�'"O�ȓnU�D��T�2L?odyB"OX����_�P��-�႗1sP���"O�}��A �dg�fH��fL�YS�"O������e�@�c��ګr7R�ї"Ol���,'[ߨ�{��!��a�2"OL���v �)JXt� �"O���4�@6_u.]�Vg'd����7"O&5���	q3�i��<�R"O�l�d��
3�|�5*���-�6"O��a,�Z���2�ȴPn��p�"O�] p��u�!�V���8[.�x�"O@�Q$K�.GE��3��SEp�A"O&,�Ǌ�(4��rĎ�72�Ht"O���ď�$r6��P�1P*\�2"O��9ٌY��U��L�+�6(���'�>/P��u�Yx���$?�IC�/:����Jڂ{\Xa�f�"D���P��xN�ȡ��ZZy�#糟�3�D)���P�2?E���B�u����Qo�
W�8@�M<�yb�5	- ��T�ԵL��������ɫo�Ju�s�B-�g��p�@àΊ��YbD�U�|�v���	�*hD��Ó�U��Iq�Ү.^� Yu��^,Yu�>�O�-�eT%�rP� $ep�=pb��?XVu�a!�)M����ecj}���VCɋ2�4+�"O��Y�߇)|�=���[�y���O.l�C�Ⱥ�@�����}r�,]�6���Un��\�,d˲�Zc�<i #Ρq�!js�O1LFv�� �_����U�f����%A����3�I�>@#���bVpI�w��"�����I�2!j�X`��0��z$i��U���"U�H(��,���'�Q���8������9X�8i���Đ�HH�c/�8LQ�O?`yhCn�1)�6���	"���	�'���g�ߐ-	N������N0(�'��L	�՗0�V���O�>})���!!����*J),@�P�n&D�( �
��Aр#Ht��i�a��@~"F�$�l����CQ���D8���=@
����O�~RC�7 01��U�u���wC]�H5����?WsJ��a�҈0�\d��%E�A(1��Jf�0�L��*��6*W&{bFI�ȓe��%�Q@ʦg�����@&̨t��L��	��EV�8�*�z���<GLTͅ�JM��JQ�3H[�M�q�Z:z�84�ȓ���"F�T���Ue�tk��ȓ0�fM��MO�VZ�l"��X�P�1�ȓ>����^:�"���L+�U�ȓj'��r AJp\N�ƫ	q�ZɅȓb h�wĜ�klhk��WtvP�ȓ
���EaĈ�G�ɽ���Lv$��J Y�ץ ���ȓ@�y#*=b��8�Rm|��ȓ%� 1�Ö:�����O KQ@�ȓa���0�AL�����[F"l�ȓq\�9eÙ�4��`�`\�(A���$G(0#P�їz��pe�Uz���ʓ3c\�'B�tЁBm�"�6B�I�~��kI�>/8�`QeP< pC�)� ���e��=FJ�!�ʹ�Q)�"O~�;$MT�fb�� ���"-��"O(v��o1�	3f.k����(�s�<��G)O����"���8(Ul�<�R	�64���K,u��[@��l�<!��#xx�kU2';�I�� n�<�5 D�T�+䏗/ �Ђ�ON�<��c�<��� F��$�d��7�B�<aSn[ J��Yb���w���Ɗ�~�<1�+L�!a��S"� I��q�`J^{�<q��ޛH�z :@'��9j�p7��w�<!$��u�v�(��F;vӒ���h�<f�L
=6�Iɵp��vEb�<y���5"g��B+]�T �`*�I�<���?&�E����H���.�n�<I&
O����c�͐z��za�f~��	�%�b�"|����-M:�U����b�<�"��,��m�FD�!��m�!Dw�{��MQ!%O���T'48����9t���p�O��[��P����Z�Ş<	�RՐ�)J���*	�'��;���{L�!(�����JPZ�C�X�#� �	?-=t�Q�醠!
N<ʖ��5f^C�I�3$ 4������"��,t� �3n��5E3�)§�X��F1{o�u�ڃT��L��&�ف&@M�K�pq��� )ʾ4��l
��'�-�"�*O|���ą�i;��`Rd")��Qq��'M��&?Ol��`�U2tVE�$�
�]��O2H�'�x�SG�ʣ#`z���F�9 �;�}R`""I��Fo������A(��q�cM�aS�c0hE7#�!�Dv�rU��E� Q9�p"m��j�P#�$G%?��kM �MSPe/�gy���RѬ}96��%0܀8�!�/�y2o�9�X�iş
"�*��߿&�v��G��dV��$�_�{���D��d���[��R�vP�"@�l�z���E �
�#K&��q!l0)�D�E�ϕZP���LWB!�DN����K���%Dj���'�HtqO���Jz�,0�L�&�-�}��R�e� ���9�p	G�@Y�<9�,JoI�-ف�n0`	4c��SM����β]�����0@�&�E�,Oʐvg��,�#���aʼ���"OpUZpa����;qLF�/����W�eזX�#X�SGd���L��ax���G��`��V��{�+L��p=��K��F!�W/Z�+Lf]j��Zh��A��LǒI�L���ȅ&�B���s�l9KӅ��-f4��
E�`���HH�.^ .$�9a�I�n�D|j5���7]�@�N�4�u��.��4%!�\���Pri� b��YA�N S�Hd����!e�"�U��2�<�EJۺR�m8�*z�bݳ��O�Ѱ�}ZB�(w��+?4 	�N�gШ�ӡ)�GJ���K�@��z
Ǔ?f�H3 g܏1���fѵ9��F"����F`���%��!3��Ux�"ϞJ�r�8��S�-�
!�*OJq#�JC����G��
��+-O�d��/]���A��L�2�D�T��**t�A���f2\cP�G��y2d�	�d���d�7� �˒�V)+��M��BޫΆ�quH�L)�O2��3�ɬx�F�J�Ɓ�V��b��^cX��d��h&J]�1�ݜQơ{�C��A�"�jI?���4m�G�D�"Z0`��ۓI�:��ǀ�?D>����e�<}��U�?����
�tJ�'H�a
���*:�P�2%m�%�WJ�Nٸ���
@�8⥛Cb>D��ʡ���q-6�a._�uO��z'Z�\�=�j�-B(b�[�HP�71"�ɧ�أ�ug��x!��U��y�H�F%����&I<#���r��0?�����?�2�R�[�Ne)�ϖ�;��1�<Ic���W�\��l���aY1|��L�(�nT8���_�B��6�_<�f���Ӭ-�<E|2B	�%����,P"y����C���EĶAd��CScQ4���I�i����mB*RT��D��)lO8āuY�8�&�c�.������7O���sn�O�!It�_�h�8ŃqA�X/��`�"�dgx�����uW�V�d��j��l��x�$$�/�y#�+_�̨�B�j?���7n��u�����m٬
Ⱦu�pP�[�6�Z/��M�;:t�Yww�lQ�6�X!3_\ܜ�k�V`�� O� �P��JL�J��dG������S.�_�DD�����i�%PX%�Q��B\�
����>IP�^q[�\B�#A�.b��9W-Dx�\@�+Q�n▴;S%�dEj4��GO� �RUh��
&��!���*���	�#M��`�b�����c(&=E9:D��e�P�&�88@��9%5P� �FM�ZFra�U,�ÇCz��1�@Ҩ)l��aD��;m�Hu�ȓΘ{p���-m�ȈGCh�H���ّG'���*���05�D_����䛳W�F�����Ru,�8��̽-��񤅣Lj�����7t���ʖ{L8ȠN��+�0�yGOX Qi(m��4O*ш3��C�N(��h�"D0�'N)��`+U"E2��x�>0�q��|=,���Ȃ;Py�ڶ�_7!�<
ĲHѡ΅,?{��e�	�Ju�'���a��
�J��D$�4]j\���i��d��YAr�+��]'鎁|W!��;�ԩ�d��tMP�ޅ]7@I��B��FNx�dC�$Eo�\�q��>	���Uf4��Գ3_��Rf�nh<�G��j�lH�A�[�,�jP�х�k��أ2��]t�����n�2�#d�*�b�e��Ն�I�Q2~y5��j�I&1"Pf�9bt��g��v�B�9�rA�	�$f��du��b���l#53��� '�'<A�8��HD��Cs�O̺��h�F�<q��%)r��8�$3�p4B��GJ>Y�&o�i��&�(��	�N���F�-�\���ܜx��B�	"�J�i�(K*+o�y!�@) �v R�D�f
����n*�O\U#�,�0[G�D�l䜸J6�'�N��Bƙ�$��dK�pRl�S�OE�.�-�c�P>s!��:h�Z`�BL�E��҇ �%x	�Oa� '�;5P�"~�f'J0�@lI�KU�7�8t��\G�<a�⇼�*օI�*��*��A9F�~��ũ1�)�� ���:�Sp�$mEμ�B�9D��C�铃I6��8��e��@�7D��RP�>=f���R%����7g7D�4�1��pNl��h�+�\uQ&)D�t��#�9`8ɂ���"v��W.4D��C ʍd�j�3���Kj
Y��$?D��#�͘*|6�� �4p���؂$?D��@Ǫ�P��еM ::+�عW <D���
Y�Um���(��v�� C%7D�D��օG %S��ސ1�h8r�4D�hP�'�3�����8L��1�,3D�hQR�A������-ԓ8�yt"6D����d߇ev,���hвV���3A5D��Qe$�//����hS�~  �k��1D�츥�ȕM2�A��C`���0D���a��L��ƍ�5���Sd0D��"�dO0Pnm��#��� b�B.D��Kb��e�҄a�b�4,�t!RV�+D�P��jL�'��c�5WR]"�C=D�h��(Q�j�����Q��.�*T	=D��P"�T$��GZ�!+Y"��9D�6�	�%��,Zv��>Y{2!2wm7D��0�W�S�ʝ���-n�X��1D�H��Ц�V���V�'h^h�B/D����,[u�4�r��.1p���I0D��c힂.��K2A�50��I�6�.D��ˑ��kh�mQ*8 �:D�ؠƄJ�&�ZQ�)z��8�K%D�0:t�="�K���|}t���d$D� �0���(!��4K\,�f%D��; �ԏ >TpG��,n�(@��""D��4�ܬI A��B��4����?D��BB�ы
�v��vI�~1Еa#D�(��j�M��d��LJ�?I��hc/-D����@�P�(���1i:��J*D�d.%��\R��o�z�#p Z�o!��M9
��@3� _hLi���<�!�� �Qj	M/E�P�S1j��4�� "O��r)�>Q4u;E���e��\�G"O�U�ׂ\�(@�1fJ]�%Hb8�"O�y�b��=j�@���V?S�U@Q"OҔ��K�Fg��8�.�7���E"O�c$H�,����׎S���	+E"O��
V"ڶQ�n��Ue��,3"O�Q�`CP���ؓ~�F�Q�)D� CG�Q4~�-S����F�$ɀ3**D����פzkT��/ƔY�L`��(D�h"��'|���{ G�D�ܺ4�$D���F�ܩS?D�4J���8Afk!D���S�X�x@g_�C��@)�(4D�`�H�]�&^�ޭ�1�&D��W�MQ�� 4N�$�
�*�$D�TꀥF@&C7i�	B�挛!� D����Hs����Q-ذS��#D�P����v�]+ccFo+Ȍ��"D�\#�k�~F�SI
?���{�n D���CŔ� #������	-l�Xd�=D����h�*pȦ��G�ef>@��m8D�xё'�9>ڴ58�߾0zԈ��)D�DІ�!Nĸ��B�_�XE�8c0�(D�\�u,��O.�LY�
�{��:D�\Ё�@� ��h�q�R!6����K�!��� /�����+6��xq,��d!��!n���H�aL�(���"*�:�!�dG�L�hP��K7���Tς>7�!�Z�SE`�32mM'k�X,��N�&}!���6m&4�t��@�tjej !l!򤟫5�bh���1� �X@*_S!�d��X��[djR�:��,!� �q
�'*�<CH�y��`#�ێ���	�'��7&�)�4�K���.3���	�'<@e��S�=�CB�)�����'��C1��D�� r�u:���'�h�S2kRF�L4�Q���
5p�'%��@�׭Y���0a`���py�'ĎP�`I��& J!+��˒y��q�'�t���k�`1���C��w켴��'e(L�R�A�m?l��1n�o^d���'�`�A1�I#>> ��FO���j
�'i��@�̀�0-,��s��/Kr�$8
�'��1i"'	�Ӑ,�S$�==�	��'���@gɩE������6J�!�'�|X��"�h��Z�%��p�
�'��[�T#!�p�ai) �"	c
�'�(�g�A�x��i���$ x>QQ
�'�rh�����+~�jE��O���	�'J�5�&T,�=[���|���;�'�Ba��	��(��E�
:l��P�'�J-�,�(<� b�,K�'Ŋ��`�
�a� ���!�o]���'"��F�˾7��sU�D�o�D<��'�B�
���(����m�ֽ	
�'��D۴S̖a�5o�4fHyY	�'.�P��f�1�D�u�U�:���(
�'����qm�4�n�	�/�C�@�B	�'�T���a��g�R<�֜@jθ��' n	��Ji�f쓶��>Eh*�J�'����SG<�z����CG�ъ�'�y*��P�(hµ�E(U�8�h\�	�'Gv�9CaY�7O*���i	�c�J�'��l0�	�P��T�b*U��	z��� V̀D+��Iy`���z����"O���t�I���1C1��p]ұҒ"O84���Zm�6��3���+��6D�1R�z&6k�n�!y���(Sd4D��g�$P� �S�aݪ˒�"��$D����L�?��O��p�`��/D��h�(�/!܀��<9�T���(D��{���j�������ꝸ�!D� B���*����
�#ذ��a3D�xq�&7$<d�Eŀ�]��Tz�k#D��aƊ�(L8�y�uAQ9$�v��SL!D��ˀ�H�r��yB��>A���&�=D�Ī�i�,=6�{�fM1z�*y��j=D��
b[.e�9�A:Z�Ӓ*7D��� ]0ǂ�"� � _�b�'D������3-F^؊�K�� ��|�b�1D�hc��� 8~I# ��EL���2D��y�A�p�~�͈�'�t�C%D��SK�U����%��M��s" .D�l�cϘ`�`#�A�	�:qh,D�\R n���,��%暐(�C'.D��r�	 ����Z-&`*Mʖ�>D��23��{�B����]5Sm8��F;D��)�Z��%P-N�b�2�"�=D��#�������o̔@.���:D��!@"	���@�z ��26�5D����Ul��8�(Q������5D�����͹v�zp�fL�0���3D�zr
j�l�qÐL
�db��1D���@f�! h�P��M�260AY��0D�D�w��b5��Z��W80Y@�"-D��JV�ڛ%w*��aC�4Apq��@&D��Y��Av�&�v \�`1Bu���9D����4j^��LS�3P\�P���0�y2m Tc.�E��#�,���f�y�ؐt\��&����5��Ň�y����j����P�3`>�)�G<�y��<oCP`��U4�Z���
�y2�:�H��,$Vt���5�y"��FV��C��J�PLu��G"�y�ձ[[v�Z�,J(G(�ȫ����y�!U�Kv��W�-�f��ե=�yҬ�����$N]�����nB�yr�N��E���n�����B��yBM6j���)�8	"���
�0�yb,�U���\�(�+Š��yBH�w�
��R�N�~��wJK<�yB�^VrY��@K��<K�'�5�yb̌�j�0�)sF2y�4��-]7�yb�gV���7i�+p�$������y2"��	@���#/��m����Bܖ�yҤA�8�HXBA`��k*�$�eÝ�y��_}3\���V��1 b�9�y2���(���
��J���A͖��y�?&4��A.knU���-�y��P��3iI�������+�yR���xV"y�ChM9 ��)2 ^��yR�G*w�B5a��!�X�a͎�y��B4n���	"cV5`d
��O��y"�I���hS��A�T�nPH�����'ў��t�cʑ�/�D����
�;Ŝ=t"O�X D��L�����+�>p���0�"O�B��ߑ~���%��i��WJW�<�%`ӭt˨iR��ԚHI2�0�#�P�<� lE�q���Bd^4�7�S�~�4�h�"O:����Q�A�� ǭ�#�:��"O�*U���|	�M �6;e"O�0�c�##Y��0/P���=3"O���3,�Q鰡�n׎%씹Ö"O i�3b�;b�"�h���'	�Āx�"OF�Y4�-8ڥ��"��]��Tp�"O�|��MԻ,���j���K�r|	�"O�� �$�f���Rpa�v	�yJu"O6Ph�h��p W�2��1�"O�!@�f�P���*�@���U"Op��#gP@}�Q���ܿ=>�+�"O�Y��]��a�7�K7X��� "O�x ��Jx��0T�R#%
�а"Op�����bD�w�҇L-K6"O�Li���
"ys��8�$�4"OF�6�ޮ=fdiq�S�;�X��1"Oč�E� � ��j��;���"Op ���8fqV�CQ�߼G�¹Sc"O��R�C� R��Cc�҄ZQ"Oa���7(1Jwd�*Sg�DI&"O$�A�#�f��H�(��,mZl "O�`K �C6S.���(�vJ
���"O��� nH�T�����DCĘ��"O>4�6G_I���U͒�J!by2�"O^yc!�V�h��1�,YuH�R�"Oj@����/�:����g<�U�"OR�sl�aN�6��-)%6��c"O��5D�N?n-��LL�>v�1w"Ox�X�dԝKgR�ȣ,��xk���"O.@�#��5D��򔌔�X��"O�pi��4�,`3��P��q�v"O.��.�u`�UIq�D�6��D��"O��bpo�|���oA.��R�"OR�i���!㴉c���a��"O�����,.���k�d�:���@�"Oڤi'�_�p��l�t���L�\)!"O0��A.�$Vu���>9D�I�"OsRŕ�o���u"�uFT�s"O>@�e"ȭ��<k梊>eִQ""O t*AG��E��)疭��!��"OP�r2�D�0ɖ��D94��h��"O0���'����C҅�Wb*A8�"O�p0G�V��gg� r}P�{�"O&@IP�Ԃm��;Dm�($w�U��"ObAg���A��q�ڰalZ"On�S�&WY`�A�מ;A\�p"O2�+���W����@ �i8D��p"OP� ��5J<V$��o�;8!Fi2"O�0�H��2L�B��*|@�d"O>�R��.#c�H�E��3�"O����zY`�����^(�q3v"O�Y�pEZ[zM�ҨE3UPP��"Ob9r���%
���	jL �U"O"��U�R9U�ʴ�D�ʕGQ8��v"O���B��5$b~x�U��2;LIc6"O�H�l�L���t@X/,��"O4��2F̕k��H�HT����	6"O<S$b�$y$�ȓd���P�|���"O����O̭]�����cNU�4D��"O6�i�`�-���D�7��,��"Olu�@�X�CF\��5��D~�u��"OZqZ�$��x$��>-N�H��"O�S��c��q�r Ea���a�"O� �#�F�0U�v��>���r"O��+e��_�	q�÷a��*""O�Hʐe�4BĶ�23nͻG���C�"O�lX���Q]�4�BG�6�\m�"O�9�Q ̷
 e�@��'	�@@�"Ot!9d&�z@	&�M�BqR�҆"O:�"�K]<�X��*��$U"O��x��+�l��Bj'"���"O���R�q�f4A�h��J���j�"O�em@�h�8����MK�XhD"O�iH��'+�䣐Ň�#>�(;�"O�!`��<\� `/V.)�L8�"O$�"�IK����WL�� �xd"O^�cW�Л�D(ag�ɜr搈I"O���5��
c'�TY1�R��Բ�"O`�%�T>��
V���3�dTz"OX��Ez�����JC)$�Ԕ�"ODXF
�G����.�!n-�|*�"O�w/\�Ylڐ���J"� v"O��hF�Z�.��#�Q"�:�"OJ��)��~qf�(��ļ�D�p"Oΰ���X?-2�z�� 7 �L0�"O���`��b�np�n��4��Hf"O�y#�'D�q;�� 8%䰁 "O ��o�KX*Hg�X<��	y�"O�ɀh@)��֭�=�rES"O���dH�ED�<�Ŭ��b|�� "O�Q��nF�o�T}zF�3w��KT"O��s���Hm��ذ'Ⱥ\c �'"OT���	��:�V���f��mF�X+r"O�l ī(UzH�ɷF��*4𙻆"O$�A�ň.����:����"O�@1pfՐE��`H�U/��aE"O���cK.q��L���`)J��d"O������
c��ya�Q7 椱e"O
a�ß����	ύ�,LT�t"O"�S$�Ϲ;�0I�׀��n��S�"O
���&J	P�!p�Q�B��:S"O"�
�ɻj��*҉�,_��]rC"O�-��ጹE�(�Hr'�K���"O68�Cݐ3^"EC�d�<�"O� �݂wJ��;f���z)�&"O����%�"o��}��D֫j�p��D"O�IG���l�v�閡_�f�]+�"O�p�	J8���`��-��M
"O��faM�j&2�� ��2���@"ONEsBƛ�'����[�"�K�"O��v͒y
h0E/�
b� �R"O�m� AF�n�Ը��X6APb�8D"O��P�Ί��T������a�"O��f��D(ڽ��g]�K�P�"O�#��+Ow���M����"Ox	b���y��� �Cv��R"O�؆HǓ~���%ɒ�Q"O���,I�#�0�ɇ�¥;�dL�"O����Gd�Q��F/h�.��"O�Q�����>�b�ꌺ`f��#"Od�k���975hl����&mI��i"Ox@b��^�zj9ZS�]�-Ψ�"OИ�sFU����A$q�*���"O��(�3<�n����ɮDz�-�y�gЖy2�Lӵ":S,~����y�ᆈ9�ҡJcR�G6�%�Bc^��$5�O�U`��x�� À���HKVTj�"O� ��+�-��b2�^Y��)S"O�8�'�� �~0�U%�B_���0"O�˓�(2Xp`�A�SPfY��"O�h��K��X��9B�C�\�)�"O�� O4pMس��%JP3�"Oj�HB�]�T�S�K�A��Q�"O$��lP�LLd�"�!�����+%"On�+tF���\I�3�I�%����UQ-E�%�^ ��+�$4���,���F�'~�t5���M&j�.D�ȓ
��bt�(�^4���\"
f�	�ȓ}�d[��ʁ(4�r�
�~,ĩ�ȓt����I�_�l�:U䋙x�����t�����[���m�Sh�wx��ȓi�P�h
>t�5�3MD�nu�ɇȓ�d�bL�:E��bF��S ���ȓ-9hpBD Z>$|�p,(�8���W!���P6�D��$�q �q�ȓ/9�e�V��'o^����V��ȓ!R��[#�0IÔ��DʤQ�&�ȓk��0(�ۺb���0Ă(lN�ȓ.��	XA�K:p*�!B�
'-����.�Du����l�P�G�@\����0 ~�p�b�<nݰ�5(�:��ȓ�4����`<����F.p@t�ȓ82�%)v��a�	���&M�蠆�z�r��A�7-�M��b�&;K�Յȓs�<�7D!FJ���qt:�ȓ��}H�΃FT���ど΄�ȓV&V�@�� �z��!�&J�V��ȓ�Bx��K5b $�����P�ȓw2"u�R+�M8F���.��G����q�D��s �+���Pb@�,����ȓo����H�{����\�
���P�lR��T1O3�+tcU�(�ąȓJ��@p'�7! ���E�.�ȓ]D	ѕ��S�N<��,'A#�Ԇ�E���#��]�*PĔ�a��<�ȓ<���*�d�	�].�h��ȓY�&����>xX����-�8�ȓI*j�� (&:��̢.p�ȓ$XL�h����H嚉�RPY�#D���
�g� ��UKE�v��!�c�>A��)C��B��(�|U(r��)��ȓw*�P�A���BQ���э|��d�ȓJ�P�p)����P�2V�|�ȓ)�0����w�T:���+{�F��ȓTx8�ѕȏ ������>MLI�ȓF�D93��0L$��O�1T�4�ȓh���+�_Ĩp��cG����A���1`�K�@�qE�>2����I�'����@ʝ�%6,��� �t��A2�'�h����΁n%>�	�kI�p�(�'̾�����=m��\��D @�*�1�'d�i	D�M	)@���%�9��y;�'t�$g�L�,��0a�&)h�0�'��@��4�|�Ċib��'ƠU
���u	5.��j�x���')��"Pج �����Q2�'�ў"~ґj��;\hcqgC�fB��f�EQ�<Y���a��r��SBٰD�MS�<q��)h/>����D���%cNL�<�A�Ǥxe,���e�'ZݜMC��K�<9ňat�Ӓc��mO<�f�E�<� Ę�#�E%��]�R����d��"Od%�'(�$֕���ߴ�큔"O|gJ�z��1P"8��c"O^�I�īc������>;�|"O:|����r�|P6)įQ6V$sG"Oi��%R$I�<�z��I ֭jC"O�ڀϊ�][��s��V�Z� �W�d4�S�ӺZ�8�� [e� ��� ��S�DC�	����`�`t�A�0��9,C��{�|����m��1�0i�,|��B�	H�|E�4���^Z��(�L��B�IT��剉�FFЉ�C#�ʓ�hO�>m�V��;7z���q�K�9 J٘4"O�uC�'��|�I���46a�"O����Bī5���%.�+��	Zr"O��$�B �9ɕ&]�j� �"O�mj�$ЦF������JÐ�:2"O��Y��>%�Żp�ٳzԨ��3"O��3f�ΈB��	
Q�9����"O�	���R:d���["+�:)��4d"O1k&�L�w�j	���� �����"O��
��g&<��gj�=�v�2�"Or�x#�,i�d<��Z�@� &"Ǒ�4�U;��#��Ƙ~C���E"O�H! �f���I�%O>��J�"O��`�ڥ`��]���۲Z���D"Oܴ@d�1<�8(��'eV�!��"O.��d@�h�<1�ۇ`��9�E"O�4`O�{m��
Ĥ���z]:�"O�I�o_XGX����Ɠv��lJ�"O^��D�� ����Z��2�("O�8��LE0��I$�}�j�C"O��R� 	q�8����� 2�\6&1D��K�g�M�����F҈(C�b!D�L��g�90��+B@�T�`3D�H*�� �0lȆ*zU ̘$%D���hN(p#�]3�[�p�0pb%D� s ��N;>�M� _ݬt�5c>D��i�� ��Dx׀�< ݖ���E?D�d�Un�	1]�-�3C��:�84�0<D�,xs	����s�T'
���wC;D���e헏)�J4���K���3�>D��٧��4%�����,�0t�*OF��'ҍd	�"�[�(b4R"O� ���U5*a����%C">@9�"O��y㇜I�؄&�@cm�Y�"ODȒ���7GM2�� �Ű����"O�(� ��l�Pm(gI�7ň���"OҥH�ȂQG9����Fɚ���"O�p��U9h�0��.�D���"O4��� �#f���K��,#JP��"O��1��LR,2d�R�Ƃ"�0��"O�	P�L$6rn13�"�w�E�"O���^�O��%괡�`���zs"OBi�QHX��jX�CA�iXrL�A"OV���<�reET:VKr��"O�@��)�3)L��4G�水x�"OH��R�ա8x<6�ǜՀ4��"OZ%��g�M��� ���.#����"OZ����CJı�-2M�n��!"O�\�1��&�^!��IȞj��ds�"O6��r@NmutM #��N�	��"OT�cOZ)�)ŨO�1N� �"O�\��D<h�J����ق@<x�P�"O� 8Y A΁<qР%�4i�4@�ѐg"O��(k܀*���áλ/���"O�<˒�(
k�p�� �2$�"O��IvFG�M�8�0 Μ�h��C"O|*�85�j՚cV 8X�U"Oֹ��&�9��}�l�s��d��"O�=r���D�(�t��R��Y B"O�����9s��R|����"O�Q� ��Ik��x�(ʅ^u����"O�u�� �.�� e���Az��6"O�=�eL�#9��Ӏ�1RҨkT"O�3�E�#F�4�I�J>��i�"O"E:�� �"	h�(	�~َıV"O�snרCj��#��8G��7"OF%�Ƅ	#���9��/b� u��"O�*�֠@D ��DܯX��	a"OnS�e�����W���T�PF"O�����SC��5���iði��"O*�1����p���*۶���"OF�z����2ni�!Y1˚Ԓ�"O�X"��_��	�q
��	S"O�l�wΓ�C(�2�o׊ ��p�"O���0kP����O����(Cf"O`i��ƂB�g���`%��"OB��������H�T�r��Ɂ"O� 1���&0$���@�e�l�	s"O��8� ��z�p0��NE�S����1"O Qa�qw������8�V��e"O ���  �f�
���L���`"O�m�V��}�)[j�>{/���"Oҥ �a
�[7D�
C� X'���"ONY�2K��rנ�rӆs@�"O����ٓx!��3I�:_`�H�"O���$ 0�����=Q��*q"O�qf�j��l�IУQR�h؂"ONQ�Iq!��J���pތ@�"OJq^	��1�#�վ���"O��I<@�9��A sE�-��"O��� N�1z��MJ6e�60U��d"OL3"H��>�9�f}s>s2"O���Ƈ[�pf�$!V$�>:?�@"O>�2P��
;��i��#F!@\ܹP"O�xRqh���&^*v�P�"O�0P�.�*f�;�a���$u�"O���]1Q�|T��"X S��H��"Or8����S�ኘY�>"f"OXa+�*&�@]��!J��8l�7"O�yC�·:� ss��?�d��"O�	�֩�i@t$(�%�%y�b��f"Oڽr�-��U�t�Pe� ^��Mzg"O���a+�Nũ�Ļ~��6"O�$0UA�:*���Ħ��fX �"O�p���J���H��"QX a�r"O�hW��;!Ȑq*���{vn�{�"O0�*��/�
�bQ�N�4�����"OV)����$,:��?
�nYY"O������P�棁(�:�2�"O℘Fj�<qv`u��4!$��H"O�<�G�/o�A���s�D�"O��+��k�9��S�!wԜ��"O�GB �e;�*U��1H�}��"O�h�b��)-��� ��S�$�d%XG"O�]�#��Y
v�ه&ɏH��U�"O�L��%��Oe
ԋl�&��a��"O�  ,�_2D( ����L�X�K�"O�]`l]�{�v�c IS�p�x��"O
�ˡχ;����B��	�,I�"O(��o�cl`�Yҡ߯G>X�9G"O���I3����C�f�(�"O�I�䥓"8<�-���$G9!F"Ov�Ҁ��$��4�,O�z�u�"O�9QE�˔5DVy�4��]\=�w"O<TFfW! 
&��������"O��hu�oTD�\�l��M'a�!�I.��<q��];<X=�E� W�!�$�p�rds刟-8V�t�%&֫v�!�ā�2=�`�`[!
p�` 7N�!��.�p���`6m;��z$n�=�!�$�;cƒ9���׸~	|,��K�!��2?R|@���X���X�@&�!(�!��>L�NT@H�� mAЄ�,{!�O�N�*H�a�٧<׈��ģ��L\!���N�Y���e�ras���l!�D�2O�V�*G�B����j�-�<<k!�D�S�X#��\�O�@�Ael�$Q�!�Ă&HD��P��Z~$U�2�� �!�$v�����/�M��·Q"{�!򄑟A1����L��)� +�5; C�	�'�0�!d�{�p����h�B�
�<Ӵ��/0J<A$K^���B�	���ǡҭK*8ce��'9C��)p� �I)�tW�Qܲ~�B�I�2�A�!7dZI+���r��B�	�xε�@a��a\l� �B�9�B�	Y�d�If)�c�"��$¶ :�B�	�=�`A`����7��[c���E�xB�I"��=XQ�X�*2�o^2,LB��9B�����Тo��x���Z33�
C�I�P~z��n�);~�UR�$/��B�)����ׇU��j��×p��B䉘F>��[@\�Xd�C�
]9z�B�	=}N4L#���)k��PD�\@K�C䉘N�<�Q�[2G���4+^�o��C�IT����&���J���'ӞC�Ɂ_`@��N.0I��Z��	&9LbC䉿4ˀ�r�`�����Ƅ`�$C�9-C�q�o�&VC4�$���/�,C�95�Rԉ��=[r(`B)�1p�B�&����AQ7B�,9gY�?�C�	7UŪ�`֬*=�$[�J�sk�C�=wT����p�D��E�ř(pTC�?%^��qvc�c��Z��E�?PC�	�L����D,��}�f���C䉌���ϊ�p!�`O�B�	��d�S�BvPb/аTT�C�I	 +���` 1J�Z�b��'�C�aq��*��5�X��7�ݠ�xC��,AK�mA�)��-��������D�>C�	)r�`t���]�C ,ÇO	C��B`��&��r@���B�ȱ6��B䉱&Ѷ���$�$z��ǈ�Hv�B�ɮf/0P��@�������7MB䉹_IHL)��T�L���b!Cڦ��C�	�-�[�	*<5��YA W B�� lRT������0d�X�n�.C䉹cn��W���}=���BK�*C��B�Tc"�]��&�s��CN'"C�ɘw���{"�U�V�j��I��B�)� �����G�f�,e3�)�Dި�(�"O�Ma6,�Pڼ���A.�p��"O���$��bm�f�֧|�;�0O�d8�	}�O�&���&�0[����cD)F��R�'�	��FTȻ�	ف1"��s	�'>��y7�u3�"������'�tl��dT6-�4H"o�>����'I��!-]�S_�%0�@�� x���+��TpƂ�%~����Eѽ=�n��ȓG���{�׽|o8dL7V$ՅȓW����u�ƙ0y~�P-��L��M�ȓxweS L�"����%�'�&M��9,�`N!^����K,-��)�ȓm��1G�W�T+� �K�x}��_tZ�(�mA,��]� *У�����	ğ`%�|r�	��qȐsw�3$�]0��:D��cfA�'[
�s�%/\Y؅00�9D��i�A�8kR݉�O�XE2��<D�HI��SO�Թk��9G. �f�;D��RD�т(F�����33����q	4D���E�"B�$Xs�ɀ�y��
1D��X�N6�YIW�\�u�ʘ�0o0�O��d�<�U ʎbe$4	���1:�	 a���</O@��d��M��V�ֹ= 2Q�%[\!���#r����f��q�~�Ip��?!�dC����7Z>jݓ%۟!�/
���[@�'p%DD`5��2�!�î%5�=���^	v3�)0G$@!�Đ�G�x�K�IW;<��}�)��n>az�����.%z E�^��M�&��<@�D>�S�O�)��ҵ�$h��lL��T5��'���` 8�\<��J��D�Z���'m�,�)\0Q��s�ܔHk�'��� ����1��&X�>v
�8�'T�YЦ�� �L#RA^� \LdX�'WPq 7��|������ ���'D�����j�X����(dD)�R�0$�b>u%�p  �Y�*�n��$��$ac(8�B�:D�T��-�(����և���T��`v� D{��Iλ}�L��"��B�A��-k��	x�l�D��`���]�$Q`�>D�D���G0i��Cu"�4D��D�<D��Ya��%�L�����R��B��9D�X�C�� 9���k'@#�]Њ:D�4�C!�&kD�E򳩖*s��cu,9��T��t"����Id��Y��S!v�|d+4D�H;��
�f��Y���%$�xX7Os������H�b�2eτت��$䁝^Q:B�Iz�(͸�l�Lm|�����!	"B�ɡ1|0xĂN !�^aC���M�B�Ɍ z(� #WV�30�+��B䉉	{��{�.̙��I�s�:1��B䉜\�}a����8`5rڱ��B�I+��[�bյ["���-To�<C�?A7���a�(k������=j C�ɝ}��:'�q��@�!��B�I.&�,*Շʏc%�%%+a�C� K�����k�+Jy��5����$5��.x=���5B��~��Y �̿ؐC�ɍ;�(Y��Z�B���K�2�C�ɮ`�,B2���/�8	0��Q���I�L��I������$räP"��I�lÆC�	�;�ؙV�� q&��Q�φ
~A�C�8<�.1�v�;c�r$�v&�:k�C�)� ���I  7"]��"ٶU���q�'<ў��A �y������>Q�b)igh?D�,������t� )^��pp#��hO�ns�{FNQmӒ�ѣG�U� ����,<O~P�b-���R���2|�2�"O�E��]3$�rd��Z�,�$��"O���D� H0]��
����("Of�
0*ܯ44����)?�����'��O�w��V������n$�ܡ�"O<�Fĉ `y�H��G&K#����I]�O�X���Jչ� ��ĉ��l@�'�B�J�l	�TP�
��#y ����'|����5Z�`3��nB8��'v����S0����vDL���'a~��*Ԝ�Ma��(h�x%��'1��!蜄7ˈa��@U��'�~�a�F3Ųh���
:I#T����d0���1���" 
8�m5�Ƒ-�!��	2W�0���P�H�"�xg$�!�d�W��$�`��3H��g��"q!��
x��Q'�iD��r#6w!��)&h\)V���RB��qq!��z�8�À�6ў�+Q�[4�!�	&T�E�ӄ+ �9���)>�!�X�*6�K�dS0p�����%}���%�O����@+X:��cJ�L
��@"OZPK�G˲Z$��`IT�Q��)�"OV�C�
5-Մͪ#��*O�h��"ObH�cԖ1�Rm;̐��"OB���� �=X��Q�c�L9�"O>9���xi>@���]�?c@u�"O����'H�XB��P�ZUB�Hg"OZyg�ƽA��:��Z�ID�`��"O>�3򍒙vZ���*">v�0�"O�<��0X�@Jqa�
6x�C�"O`�����'�u���X�0.���"O�49��-Qo��!Ѧ�$H<�9�"OZ	b0�@2	d�#w�#s�h G"O�Ԋ$hǣr���k��^�VDU��"O�x�ۚ^˂��\�"�"OHM�S	B48W\�Pt���!��tP�"OZ��r��'���a�a����"O��׊ί{u"l�u �|(���"O(��Θ�M��z����j]�f"Ov��tK8�ce��I�TQb�"O�u.�3��o��+?gz(*4"O4`�'H܈!3.P�H��q�w"Oz�g�X? Y0U�e͊8b��b�"Otm�@��=%�����l�`"OTBk��Kt�H��Jؐ~|؋b"O�����F
z`��OZ�v����;<ى��Ӭ�����/�@i���d��m
DC��:aG�E@ �'E
��S掌�C�)'�"� 5J �q��(�`J��&C�	B8�u���Ʀ&zܜ���Q�b�<��F_RN��:�H�|��52���v��G{��-8NAلG��Hh	� ��y�B�(�T&�1^H������yR�'m�'3�)�'u�ͪ�h@�pؐ��B��4M�ȓ��xb�ָ@o�L��M�@�Tp�ȓ�&�c���h�`� ˎI?���ȓ5t���R.Q>>Ե�"A�S0�ȓc�l�MGn������	'BpFx�W��D�I�#Ot.V�q��ѻa�#�y
� �mc�B�;-R��F��I7�2���O�b>i 4�\,d��qDF�7`X$C�+D�d9T�H�xi(���_0k��\��"&D�l��U�qRN��C�+�h$D�H�'�4�b�2Kf�`����=D���FP[���ױ?�Z
�G<�I꟬�?�|�����Q N)���H&c ZYz� �t�<�祃�b�T�1f&+;4��%�Ng��?�����F'#S����U>#���Q+��y�E�Q��:�DT��X�U@M��y���;V }���
������I8�y�h�{�֔�!��"Ȳ��*�yRɔ�^�p������PQئo�՘'�r��iJ���ț�X
�ۺosPʓ��S��y�Ģ>�d�2t��x�����*V���'�ўb>uA�JI�-^d�����F$z�h$D�\C��@����	�B�FB��G�!D���]!A��5�REخ���@�$D�d1s�;���Xƀ� 2���c!�^�f;@���X'D�v8�t�ߜ<��LG{ʟ8uc�dD�uJ,��c����*�8O��=E�4/ɬ|L�i�a�]�)|���W�2�y"�A�
.XP���B6Ơ��b͑��yr�-��uе�ĩG��䁃Ɇ=�y"Iǭ�X��Ä�G�z]��F��y� �V��i3�'pgn,PR�զ�yB���O�֘�a�I(f*�r"���y�/�����h�΅�W���D*�yr�׷K�&IS���y��x�Eɮ�yBg�7^�Z4⑋A��Q�ыV�y��
7 b:@ ����1cQ�ɯ�y2� 45	�x���*�mף�y&E��^l�P�E 
�X33��y�J�D1��� zJ.+TkG;ވO��$�O��?Q2S 'QJ�}� H�JD�Y3`5D�D��A�NK�=`b��F��0�o/D��h "�wFh�P�שL����,D�ёb�*�� ����)� ��5�5D�t�D)ż<�R�j��.. mx� /D����k�D���[�+�V4�*D�|��ɫ6�����Y�u�إ�4%"O~�d�O��O"�x�I
q �aP��^�q����"O�"oU�����K.��"O����_��"`2'|��=X�"O�]�W�^�{a��Y����RY�"O�Q�Ԡ�%�����d�=*p��C"O�S���X��jpI�"O�P�Ё�;/�FxF� 2����Iן$�	M��/�F�Pf�DzT�!�a��>4]0E���y�.A
ph�?D��xDH?:��$	3LA�2g�@��H9D��@
VCdlI0O�	)��㵊:D��)dͨj������,D�z�SN9D�X�&c�u�ibڎ禐�57D�t�T�R�dc�W�M�@���3D�l"�GN-3K6LҌT�O�85"��1D�4���ϵL��,"��P��� �@��W�����_�]ٸe+VL�/G	l�9D�:K{!򄝃����J<����`�ўx�!�d�`�����P�����C�s�!�DȍC�΅���^�z>�$�#iЉq�!�W�Ec��1fשO'����żTi!�$ߕQ��5c�kȺ;~B������W����݈��� ��}!s.Y�|�6���"O� R�A����Q��d*�8co�c�"OTME����Ta���ZՋ "OD�aA�W5r���� H|Ɯ�{D"O+�+�<2S:�� "Z%���[�"O�Y�B����1BP�9��	�"O�I8��]�{�4������8|��"O���%�:�D���o�X�	IQ"O��sG@� 9�x�!OP�%O��S"O>���IL;�H ���1JD:�2�"O�di7 �.G��p�-�&b`�"OD˅�>��|�녾ENIj�"O$�Y]��]�iP9[<�A�H��yHTp�5��</�l�ag_�ȈO6�=���K;��¢49���W/b!��<����	ܮd+����"=�< ����Xm!��P.4� �e�#$"X@U��W!�D 'P6ȩ#�ۉW<�*%J$/!� I��|G�5*����1"](!��E�uC(�	���~�YrAҸ7.ax"�	�Y�0�{b%M�]:�er�r	�B�	 
x��C����#��͚V���c�F���6ڜ��.C4�����6=@�A�ȓ28���b�;J�j�Ӄ��� ���.(J�*ɠX�V@���F� �ȓ*�Z�ц���z�z�RG[-9�J0���u�RN^�;Y:@�F�Y)c0� G|������ЀLɫz�=�tmT?�bC�I�/s$T�u�r��@���#}dB�I)`�d̘Q��� �np@�(_@��ƓY.���ǖ�N���$6��h�ȓw�n��&É"�l��d%D=q�фȓv�J`IDY*����M�W2���N����A�8'%�0� �5����5���Bw������j��H󴬇�`y�02F�U�l�t�R��Y�.��P+��?�1��-_ĬXq'��t���Tj ���x���G��R��?Y�p@FA��y��V $�i�vA ����T�Ȣ�yRO	�;�&����A+(����6�� �yRa�M��d�LE�$�w �5�y�B=+��3M�7�
��Q���yB���H�>1��z7��aT���y�h0'(��F�b$�S���yb���������6�q�M�:�y��ͥ���q����R����]��y��FYb�ፔ�30$yWK̅�ybB��&(
]q#� )"���Ʈ�#�y�3����&Ee� a�K�yB��SjD�z��Ȳ~D=�шԑ��#�S�O�QY��ĝ��<3��[�ki���'b�`�r��XZ�\�!��g6�X��|��'����yZz qt��v9�93o��F �ȓp����3Ǟ�]�2��U�~>@���-���"G.@�yb�M�e- C�a��D2B�i�l��8҅���  s,BY�ȓ@ Z��RK
 �dPr7G��x�D��ȓ|u��y�ǔ
%I*�8�Œ�3*�����dK��y�Ha��
�O(h�L>I(O1�1O0pH��ڦ9�а[DQ��"O���)ıF� �R�O�AS���V"O�mP�֙:���a`� �DЙ�`"O�ARE�ֆ�����g� ��S�<��F�{*�AJ��;1grЛe�M�<ѧ����XK&k��p�s͝G�<� Fт�喺ni|��oO��|�V�%���O����� ��13�j@;�&=�7mU&�!�ŌҤ��8A5��
[�!�ɩk�|����ɭfz�e)A��&�!��F��`����G�����.7x!�DŞ�x� ��H0�֕�G�G�!���7"�8��D"����q���{!��7S`�$c۸l����\�.h!��@�֤ȧ#�dZ�݉2"�2X!�]�6OD�`a��4Pf�G�\/=D!�$�u��("��ŧ0?H�4GA�V1!�K�)s\k�f�*?lEC5	=?"!�D�?�pLY��f<��#R(!!�dU�g����+�����S���2sn!�D?B�:|Jf�C�$�ܭ"7b�
}!�M<�|��RΑ�d|���̘-�!�$�lJd�%֙9U��!�P�!�d�$,b�$���C?Z	#bFT�!�ަ@��eY�`��u�Vp���B�!�d q�v�@KJ�Y���d� 0�!�$ύau���o��Iq�24�59'!�d˥,��t��1}aP�9ģ�6%!��	��8'��C|e�'�٦M!�Č�-_v���*F-KN�@��-��%!���Lu���>`�<���G:j�!�$>?{�p�bܺV����/p�C��$�`(�w
R2hx!�т�>2��	E��cx�@{��%Xj]�v$RW�U��7D���[;���2I�
pӜ!��?D���bf
�PAj#'��DƈM���(D���סU���A+��w-��X!,D��3��Ɛ`F,�"�_>mp��J%D�xq�a֍O6E	�]-,�ٻ@�#D�,
B�[(Ԭd�i�S��t�҈ D�,�#�;-���E� ؔQ�" D����NQ�U�2�¾>fdZ�:D�t`/i�]hˀ�s�4�֨%D���'��_��1+#�1{��n#D��paiF��@�@��b@O"D��
`eK�64" A�c]CW���a� D�l��F!Gx.i���ůo�K��C�ɻ9����p��*364Y'	�! XB䉖~��Œ U�nH�C�U5��B�I�[�#:{�1� �+6i�C�I-S�l=�M�i�)�󯆗RJC�	�|�#�cƺ%��E��D>�6C䉾B#Z9�ԅ�"��5���t&C�Iܸ�J`�I�(5���gM�4QQ(B�I1R"��p@�R7m�W$B!`E�C�ɸ0�l�j7��'%J�[��D C�2mr�` �ݾW!H�` �R� m�B�	&�Z�� D�T����t"ۘq|B�I5S�v�1B�� m���rB��B�	�*Th�R'��32�٘5��!��B�	/rD��IE: @P�a��$aAC�	��Z����|��:��V*vC��{������Q�y���;$C�I;R�@����6;�u0C�R�6s.C䉋Yhb���$x8V\2rO�D�B�I�^1 �0bJ��pN$(�J��[��c��D{��D*�s��r7/Ч���	���y��JN�Ji�@ɗ�g��X��
�y��f�����H�Y���
aG��y�B�;�rXW![=) r��Q���y
� �B��ζE��� ���H���#"O�)@g�"f����������"O�cAP� �Y�SL_KJ���	x����@\@���K(Qx�HS��VMh<���>Ĵ�P�;=D��k��l�<a� �+v�"Ao��0�����o�A�<�g�L;.#r�{p�
/ �0�80mAT�<Q�K�?2(��&Ȅ0;}L��(�E�<qFKZ�XqI" �{j��(��<)��² =f�:�]^�!p�뜼�?ъ��9O4���rR��1$Q:�23=O��d�2h�~��v�R&�`D�#��<�!��s����Ij��!���0�!��rє����C�Ig ��fe�e�!�ę9���۱K�u�쑱����aZ!�G5HG���6���q �eY!�$�(��L	T�ɜ�~�bc���t!���Oi v	�!т��2N&C�`��u"OIi���	�-֦k؝+�"O�
r���*�^�e:	r�"O�D�p˔3��b�Ʌ=a�Hi�"O���Ӧzs�h��h>�5"Op�`tËV_���  ��g"OvPSWᎴ/�f�q�O;zp�s�',�I��r�ؠ�&�hb�	�\�@B�+x�萵'D*q��ܢ��?��B�=��b<F�С�񨆟QtB�I� �t��v+LWS��#F4(C:B�I?�H<�&�W�k��ИD��x�0B�I�+W ��K�̙�ɂ5ҼB䉘x�p8:��k�f�M�2�d���=y�_2n�i�(�m$X�0m�0m0(�D|��S"����ŉXQ���0� 5B�ip�2��QϤL۔oN��.B䉔x���Vg��_�6��U�
"[®C�;d0�p3sG�p�A(qLD�(lB������F�jL�*�B9!�fB䉟n|��j:.�b���x�8��?9ߓl �إ!�M�<]�����XM��XEA&�L;zR@�G�=��}�ȓa��,��7|�0A(R�ҜE%��ȓq�6���#.Rx0��_�#v�M��4,�pf����6I�@��*<z9��2R���-�1��J�K&r��H��R�:�fܽ9!�IrAȥyؘ���Mv��1���<w����D"[���'���'yɧ�@�Ӳ�S�L]f� vHDL��%��"OB1�#G�0$,��(V�]���&"ON��q��k�$dѳ�қtL4D@"O�	�PYKJ���aL�[<*!��"OƉy���c, �c��*�) "O9y��.K�b� "B�"k:�P"O�e����'�8< �Ǖ�T��(!9O��=E�dH^D>�:��M�@A�P����y2��3 �l�kVʁ�	����
˷�yR�G9h
D�$)�,��2U#�y"�:9�(���-��*ʝy!�=�y���'�8\+s��, OP�3v��y"��3rD���J	([H��@�4�y��� R4�4�ИIm�,�6��y��N9A��X8��G��<�H��^��y"fBK� m��c{N���g�
 �!����(`�m��ȡk�EO6:�!�d��ocL0aq���0� H8�d�!�� `�)q���kÊ˲\3Ab<�"O$@e�ֲPM~a�#�g;���"O<x��B�R#���B�M-�A�'"Ol4�4h@)@7�)�'�O�*0�KU"O\Q��o�2~:L0���G��:@"O�T�@K�v�L�Q�$�80� {�"O�1t>x���3�����=��"O}k��kX��a3h�Ypd"O����E6,�80�"[D!�"OnPa�҃~: �K���6)���#��4�S�'D�z%�f%��4e�a$ڄx�����B�v8��<)J�ZDިaz5�ȓ/�Y�i�$�������~������.Ʊ{���2b�C�7�@���y��֋��D�����I@�V����D��P�&�	�~- W�ƪ^����ȓ9'�I��BN�( �n-W���Gx��)Ea��Zl� [�|J��F�
w�<9U@IE��C�L��vp%�y�<�S�)�8����2��"n�p�<1�N,ܶ܂V�O� �����m�<�F�	�4^����/�-)=^�� �R�<y��ȡ��e��$OF�d�OS�<�����Xҵ�A�����Ɗv�'�ў�/�<D��̔�g�lH4$E�5��`��pw��ь�k#�Üh%���Օ!�ͿJ�蝂#���
P���"ORYCt��i h�hQ�%2��[�"O\�BF��^�jq�sh�g�$u��"Oܰ�""Z�W�B@b�G	.�x=Ru"O�qq�=Iy<�gR;�(y��"O��{C��0{@��&�H�$x���"OX���h����X"��B���1"Oj� �
UC��F�,h���R"O�-��擻w{ZH�4�*Z�9�"O>�3��R�p)ڇ"�>@���"Ou�A�5�
X��.G.-���"O�TJ��^�I�RE��n�qp�]C�"O%H���-nZ⌻0.�,GVYJ�"O�-� I�J����2��$J\�53%"O��ٖg�6�E���M�8��"O�ћg�(��X[��X�l� #"OډxTH^�_���`���&^���S"O8��Qd�(&d�P�kF>$^�t��4O��=E����JX���q��������������>�S�O��:R�E�|��u�Q"�&K�݋�'wJ��a�[��>Y С�(?�t�8�'�6�Q�����x@�B�%��y�'n�y��'��sX�()�dY	g�tdj�'�|qQ�ٙ	���c�6a�$hH�'_�}B���8�D��l�R���b	���d܊;�"a���|���V?8!��G.-�h�ǀH�<XB(L6%�!��6wL�T)Ï!2����@�(!��Y*�'$���(��!򄗝4��`���?3l���H��!�T�C6E��M-��AI���[!�[�}���� �X-p�f�[@	�4H�a|B�|��,R����'�h�Tl;���y&��?��ǖh�&I#�W��y���#�px��k�0�⥐��6�yr�B;~* ��ci�7$I���g��6�y�A��c!(�� �S�M��9�GШ�y���*��0@��ED�-9�S!�y
� Ԉ��/t���L5h�L1B �'��	�A��{�Y�����b�Dz��C��vd�4�V%ڼ0��ujeE�(��C�ɹJn�M����j|�9���K�bC�	a�<��A:)�!b1�%�2C�ɵI	
0��ۑ;~�@�嘋5�C�7Yؘ��m��@�@A���/6WC�	�Lb>�0�  _hތ['K�=��C�=A���$��i��Lӷ�@�G'�B䉁Z%xAV� �P��h�$I� E�B�IHrHI��1bMi`�0ZpB��!�x��� �e�8}�Pj�]��C�	B�T�3�&
�sm��aa)	���B�	-Gl���t�ٍ����b0z�B��k.�y����yv'�S�^"<щ��?AF
�c�eЖ�\6$&��gF0D�Xi3N*PPH����Y�$�ȍ$I D�P�%mJ7hbP��g�L$�qs�j+D�Q�>�pY��L TK��$D�d�����"�(� `���a�$D����'��1ѕ��EX��;��&D�����fA�a�6*��|���#�����c�͔E<(�4��-E�Q�c"O��&&�p���I��A-����"O���irE���#�\�Y�����"O<Q��	5�=�����d��"O��@`��(C,P+�l�#�x1�u"OJ`����1�H�O�2���1�"O�a�4O
 ){���wDm҃"O�A��9��ء	�6a��DZ"O\�;�BP%[>��Ó�J+#��"On%W#L�A� ����"XU�"O�����=�ty��ϏEy�0"On�z��4ey�i6m��5�b�@�"O��C!��r�Q����zˈ���"O"�bc�X�R�(�˅�wZ�B"Ot@8�/G,b�5kS䂳eY�Xʐ"O֐�'���U�b��4�ԎD�<I��i�(��a�,�� ��g�<y<0�xx�E�]�\X�cHd�<�5,ڶ3�2&盆��ix4�z�<����^l���߁]M�a�B�Im�<y�.A�@��y���(]_x��#M�h�<�A嗾t/�ظE�^���uȟ]�<ё ˤFX����s�ؽ���Z�<�7A(!?�|v�+X����k�<�woW#	t�1�b�� ��HS0,�d�<a�$ȟ{��!*9)�� �{�<�p���f�*9���8:��A0A��M�<y2�ն�	)%H�5|�z�crk�U�<���
+|��D�ִg"Ja;3g�P�<�%/)K�Z��s�L��3U'�e�<1��= �D�I�Z�
��&��W�<!��ݻJ���@T�g��$3��T�<!���J)�&P16J���b�Q�<��3����ɽhH����HQ�<q�.�*D�f&�O�qf/�G�<q&�d�I˖I�d_0�/��<9I>Y+O1���q�8d80��\ ��� �&Hm�C�ɋz����&A��ά4t�C�	UX��ũ�`�(³�qޚ �ȓPj5��,�<ݘ)[�<.ܵ�ȓ^�l���E�Q����d*�|��.N�*�M�o�fp7�#{����S�? lТံ�|�:4�F"q���!g�<IH>E��'/nY*q�1s����u�Z�Q"d��'��7.FqR2��w���{�'1\-�农"���b��B�#�~$
�'����>u^@ Ĉ�r���'� @�U���%�kרߜ?b�K�'���R.�2��ֈ%B�f��'pu+������;�IJ.�
���'FD��B?Q�>�v*O<-@T��	�'~����
�>��F�E%-C҄*	�'*�[��Ƌ�6�k�	M%+/��	�'�f�c�������/*�|��'Y��9�@(/>4"&��$�>�'�G�E�t��a:�Fܶ�8�
�'����ԏ�	��X�Q��6��	�'g
-)�n\$tl�����HtT�	�'��8�^Q�8I&�ӟoI����'W�4KQ�ǁ�-�f�����'�r]��lLG��M��:i���'�
�9S�;gLМ%��%|�U��'7b�)%�J�����Qm<�m��'�L���'&6=�D�hR�gP�0�
�''ܱ�dM�_40���@\�,�	�'�LE� �SV���2P�h�j]��'d�A�b�P=I؍ˀ!��k�� Q�''�=S���"9$��
�ޣd��<��'��z,��s�jRG��
d��p�	�'PL1�T%mDڦ���0@t��'�>�z��D4���.W�}.@��'�\�s��ܕ���c挜�n�d��'�~�NHV��J�ʂ#�e��'�ʅ7o�a��b��O��F���'NZM�e��HD�Y��)сw��=	
�'mb�#���d�������?X���
�'\z��hJ���ł�ƙ�6 P�
�'z*�2CO"8N ����e��H�
�'ڌW�)����	Ps��8�
�'4D��Y'w-1�a&��d��J	�'���FGݜ%�l���G-Z?����'8L�
Qć
�,-2Ć�W��{�'� ܛ&O�d���ѥQHzhB�'h4���B�y�sC�La����'q*ܙ�m�#�"X���5BƔ@��'��l{�iS  �HI0��7\���'sb0K���#obe��@�6�%�'����j��-��7"�C�
I:�'mT�j��Cc_bE�q�F�R}�"�'l��x�U�N�2 ���LK&d��
�'2ƴb�B��A���aOѥ��R�'���"R��BV����>�"��'�y�E��"+�1�V�Ĵ$�h��';�
uƇd'��[� M�'� Z���Y���I�B=����	�'��m�˒�i����)��䔩�'���i jK�0�z �EM
�����-D�`ɅN{6H���?'�(�+�#)D�8���9I!b�ĳ?�C�k,D���R�ݎp�������;H�ĩ�g�&D�����J |u�$j#�R!;�7D�`�!�:r�\�a�oT0}$:m�T�/D��k��ɿ9Ĭh��S4�0U�7�;D� KW��U��#�Ö�*�Vn:D� Q��Б��P[���:�`���9D������!*Ar A��3	S|�B�+D�� *��R��}6|k�T�;6 H0"Oj9��e�CO��t���w�kb"O�u À�g ��裪�5^���f"O�k� !8j���2Ĉ�3nY�"O<u�F����g�F12��R7"O���FN�!3��k�*<2$0W"O�We�!{��U+B9g�陰"O���T&�H"Xt[1��T�
Ű�"O�{5�ѳy�R�����x���a�"Ov�1U�B��|��#c�^�d�1"O\�yGlQ')�T�ᜥ���w"O~�w�ӿA���B�j҇�Eu"O~}Z�*c�Ҹ�<$��Lc�"O�=6��~�μ8�F�`�tP�"O�X�$[0,|@tR�%�6-�l��"OĭX��u���L�/�~L�"O��7��"-�fC�B��h��"O|���^�<6��J�ˑ0PTQ�"OxTꑆ��z>]�RKN�
�h\��"ODܓ�G�M����/�3i�B��R"O�mCG�1\vp82,� �Z��B"O������/��t�k��K� ��"O0`�S4�ɣ@�"�@���"O�4@O�W&�:CA<91"O6isWa� ����@O�0����"Oe�S��.�\�.��$����"Or��/֧J�	�4�fݞ�A�"O�Ib���VX��FE�����5"O���cңB� �(�� ���b�"O�ǋ\<���,�\��9� "O�%��O_A�Ua��^!Vx%�!"Oti�󀖖2o�����ױ,��"O�qa�W#'�y�&�<m"�d"O�I�*�(}�UV�8д�96"O�je���s�zᠦ�ɘ*��a�"O��胋�I�H(QE$���zԲ�"O0<(��ՑhH��sCHj���X�"O�;㇍�~��	&ᇉ\����t"O�m�`d��dU���#�֋�.��`"O��jЧ�&;^@�2D�(y���9�"O�塥N��7g싢���C�� ��"O(�+g O�5Y����ӯX��X"�"O65�`䊮3�h�CŠ �fH�"O�J�&^�Z0�2R�E(�"���"O,ɒ+A6B��S!c�
�M{F"O USGeșjG	����f�"O����	3	!0��o=�l�xU"O�E�$IoT��[,\�:s"O@�v�T;<�V���	X�*�"O��@S��7]º9�d΂�b$�i�"O�ŀ�g�+�,�p/7Y���"O�T�dۢ.�xD7�L�4Z.tXb"OD�cr)6L�H�r��
n���"O�mi�+R�z�H�S ���x\&�0"O�(�8t��tj�KPv��a�"O,�v�@�&l���ܤz���`"ON��QL��qߪ$Csh^�\ψ�
S"Op�qFɶ4 ���fԫ{,�p� "O�����+j��
wk�x	�	"r"OB8Ȑ���l#��@B�@4Z	���a"Oyڷ��++�|E����>.K�(�4"O���0-�nb��ӰB-ZHI�"O�좥 ��#�5;�c$m{6�s"O��Qw	�	�p"���"sz�9�"O� ��
�(5/���a�� `N�6"O&Ń�L�>{9����A@�iV�в"O��	�n��~%�U[��G�%2��z"O~,R JD�����o�=C�|�"O|��ׯ'
Q�%�"��9bTMq�"O�sB�ǟ#i|�C����1r�"O�\����L�ƅ���z�(�"O��9Q��obH�`�q0��qB"OH��5�\�;�t�5�A �l5��"Oh �Z��y�����3~L!�d��(1"�%�1n�Q$� pQ!�$R1 �Y"�^%;ð�d��{�!�	'14���3IR�M��ܰ���'`�!���6{��CTIң)����Ӗ5!�$�@�T�4��S���cb�4�!�dǨl�`�2rK܉&�ݸ1���!�Z"���HW�+ܕ�$�P�5�!�m�� HA�w���YЂ�,a�!򤈾�d���G20��P�CG3[�!�$�W��ur����\��}��D��5�!򄋅t��$���2^a
��/!�D���<��+�*�ր�qn@'O !���m(��'�ЎZ��٪��Q .!��9x����!�r>.�`씗v(!�D�-��E�!�+�1R��R>�!�������mT�ܴ��)��|�!�D�d�py�(�B� ��4H�:�!�3Ld h�Ù�e�Pm�-Kv!�V>�pzs��w:py�i��!��_�,��`y�F�Hc��s0jW�!�D����$��&VR#��E&M�!�d�h��`�7�4)O�9�Mѽ"�!�D֘�F*�?G��f�)o���ޢ*�Ƶx��V.�E���τ�y2͞�`Hrq�LΎf̅k%�Y��y��64���C���P��%�̑�y��L1@���6O���PS�n՛�y�Z29�y��glp48�/���yBi�:���bO�Q���R����y���"��H���1x����õ�y�,j�<a4��ov$H4� �yҋK�1`8�*f�ˋc�0D)��σ�y� '��q���UH�@���
��y�B�q����4��ESp	"����yr��R�R�𳄚�9]P����y���%(��U�׌ߘ*�b�iW*���yR�$OJ�����!
u�V&��y���:�00Յ�!Q�	��iA��y#3����+�7R4ɫT�<�y҇)Y�%3.D%׼I���y2�_!="h���줔�B%�&�y"A�yu�]H�ş���(��ʃ�y���2e�Ar㨙�1Jl{Ђü�y�#�/B���&л%��q[p"��y	܏Wn�z!ܲ�8E�g��yB΃w�Z$��f�;)D��g6�y��hnx��!X�&l���X?�yB��2'��Z��#~}<	�d��y�=�L	�ե��?1�M���P�y"I���b=��W=6�ht�'@H�y�l*n9�Tn�>+dQ�$*S?�y"��Q+f D�%�z�����y�F� 3z�x�L!F��La�A)�yb�PQ ��e;S�|�iP�-�y
� 6�Ea[)_Pt�3��W�:�.hB"O,�j��Ʋc@L��'I�Z�^�83"O��WL��3�D8�Q�)�x�3�"O�m	%�ڹK�`�J%�\�5��As�"O�0��a#|پ�U.1π�r�"O��xoND0@����zӘ��"O�8"��:Zt�,C>�V݃'"Ov�B>h`��KK�2�~iڂ"O �K A�)��9��M�p��"O^ a�ゑEd��(F��@�F"OR�E�M�t�L, FO7�8`��"O�ء&HC6K���+�k%A�2���"O8��׈	�L�bkܠy�.���"O"�h�Z�3̊}Q�D��a�bE 3"O�[CnΆEЈ��ƩſH�.���"O:�#e(�=Y��l �H�*����"O��RAP�(S֠��ǀ�K�Zps�"O�5����\����Հ-m7��h"O&`B��Y�/� �Q�K�X�p�H�"On������4� T��lm��U"OT� �ΰ2 ��a��2?h����"O	�S�=b���5�X9`ks"OP �#��&.��M1�M1_P���"OD�0 I�%o0���� �c��B"O~�	��&����[/#/`�RV"O� ��_�]}8z/L F"�P)T"O�D9RnިP�ZxҴ@
1mh��ѥ"O�M�����/� BB�K�"O�����ܢ2�4��]-6LE8�"O����o��iqSAF�<"y�0"O�=R7O��?T�����2&T�"�"O���^VW��mݼ�lPHd"O*Y��kK#n���쐣�@t�E"Oj�0��Ο�����H�m9rIC7"OeD��_B�* �P�3�tiz�"O"8Hd ;]&T0G�&h�D�B"O�岣h�p�;P�<I���"OƱX�䊅v�	�IU�]�a��"O�(�WkG�[O�L���	�x� ("O�H[�k��U�V�ꁩ̌V��us�"Oa��ǡu�p�I�3)�Q1"Ob 8�$MT�]��YT��"O�e@�c8K�|l�V��
69'�!�䇩q�̅bWI	�8�T �K�T!���=;���i�4-2����	E�U�!�ӄ{ �5���Q�4�F�ǉ\�!��ڑl̲������ǃ��!�D���^ [�
�� Y�+�.�!�׆QVhaH0�M,9&�����',�!�TK�0���V$6O��"�71�!�䜽t�l��-K;:9��*RW)o�!��v�tAW�M�O b�1�/�8�!�dA�/�Ȉ8r� ��:ѐg�(@4!�!]^N�AdFʟV��)�R-E�(R!�4k蕃��9�b�j3Ǉ*)T!�˛ r�B�*X�}_���P�R+@!��?5��ءb�%IL'�K�49!��S$5[ Ii��G'j#dU��$��7-!�DD�:�2l�e
��s�*T�%9!�Ĉ'� t�&Ӌ$)r�c�4!�C9)
��;.�D"͐z�!�$#f(���RL�$�!�dX8�:�B����9�$!��	GR�!���=נؑL�9@�����V l�!�� ��p�D�$:
�y��7"�Ʊ�"Oʽ(��B�bO���h�}�"�q�"O�� &�2��(beN�-�rѲ���Ox��*-�(p�.ȑ��Bd�<���%D��0�B�/�`99a�@���� �5D�@B��P�j@ۖ�(z����&5D�,�燊�:0+ �Cʰ)�d5D�J��Ѽ/���``P"k�� �b�7D�`��Ë9?qR��Q@�%>a����9D�l"b*
:	�:�$ȋ+Q�=zv�8D�|�D��7��96�
�\����B7O.�=�U�6$�h��-P�G����/r�<q !0�Ұ@���*X`:��B~��)§.�pmG.G�X��ꅇXl\��f��w��$�Tq휘b�I�<Y�_��@��Ŭ*����J�	���ȓj��7�L��Ƞ������ȓ����3�ф�~���n�bQ�ȓr�6��(��p�"3ZU�E�ȓ	F���E*�O h����2k`��D{��O�j�B���<(��F�A$^�nXY	�'a�Ib�@Ӊ)3�(�L�U�5�p�)��<��"l�����aP�BS&�jg"�E�<iP��q�Ĉ���֝;��Mb0.�ß��'�a|���,��}��b�̛�)�y�ƇF��a��ҽX�x)S/� �y��Z�L!ֽ;sL�Uڰ4r��U��5MQ��?�ʀ邾o� ���>n�!�2D���t�5BRH���=z�2ő��$���<�u�/0hx���C��y�t2�o�C�<��`]3Z��(�FT84�.��d�Rz�<�� ��"��0 Q�R�`�< �'Ν}�<q��+z�2����T9Rk�!Zr]v�<�uLJ ~�Dɔɞl��p��n�<���	x�艔�~�q+D��i�<��6 �<g'K&����h�IN�Ё�Y�r�&p;�O�=i����3D��c@n��]}�!SƊ\X�b��0D��H�i�Fl���G��^ܓ'�)򓋨��<�dCц>$x��1-�ո"O�h��35��� ���T����pQ��F{��)\�=�v\K�`��yh%�y!�	7��zD#E�8�T�`�%e�!��5WyX��r�I�B�d<�2�(J�!�dA���0�U��8�LXj7,��HI!��ϳ{�};E��� ��b�V�w!�1�i�WhA;���`-A<�!�d�As~���a9�h\�����!��ԽH.�īD�	1Ctu��
��!�M9��	�7l��
U��0���,�!��Ģ�v`�1�	�7Q,��QIخ8�!�d�^�0�6,�Z��#v��	/�!�ā%�z����%\M��K`�$w�!�D�$%̊LJbH��Z���H��u�!�dE2fnDYw��j���d̃��Y"i�R���F�3�$aC�,��y��/1Ex���$"�0�����y�@'O@Dh�������E��y��%=1J���.u��`�y2��`qï_o�b�S%G�gN���/��4����2�Y+�K�8`��t��A ��vf���*s6b+dy�ȓ�n����Q�y>�:5��&~)��ȓA
� 1Ag�jVȨ�$C�th����S�? ��e��#��8�MR�|�(ab"O�쨖�MG4�A��)��٠�"O~�)qJQ�)����3��3@�r�I"O����*z ����Fh���t"O�I��U i?d\��j��z2> i�"O��U���	�@�$R
�2"O�@!�b��N1
�� �K稐�"OР{e[�>h�{�m<88��"O��*�.D�j���/ZZ(��k"O��84i��"��{D�N��Z��g"Oj8X�C��0�TlxF�^����1"O�mZn
�g|�I����OHꐛ#"OL��&V�t�h\b�Q1SV��h�"O���S��K�D���L�C�)i�"O"�Y���
:dp�b��rҒ�i"O��J0fF-ZF�{�ᛤz�d�D"O��H�OP)��LЁ�I�&��		�"ODȄe�rL����/ �,�:P"O�M���M:M"\��Wo��5�8[�"O�@�F'�� N� ���"O��d��!>'M�1�ڭ4�$���"OȄ�AЫGt�U�e]ؘ��"O�9�ؾjL��8�7�"0e"O����I����
�FY�E�"O�(���Y�u�T�:���P�"O
`˦���L�	I��"az�К�"Op�@���U���ǫ� f^��"O�AE�qQzq�b��.Dv�DPB"O*(3@nH�tW>�R�	�H��T�"O�D"����f�"�z�N�v�n)��"O����N.�@E��45�n�2"Op Z&�.��8� �C�_�Z�b"O4��`�< ��%�q��f�<���"O՛7aX�`�\�&��A���+�"Oص�/�0����V&�s�B$��"OF12���U�I���f�&���"O0��Q�I-,E܌rE�OѾl�"Oh��d́�/�-�dT�q_��"O�t  �֊��I��JR�"O��鷤M�y����4B.dzp"O؀H�E9K�&B�ܐ�"O�՘�ɏ;~˨��D�A�S;�YQ"O�MQuNw���7D#X2�hq7"Oa���_( hd+��6��"O�e��"�)`#�)a�! ��`��"O����Kf*��G`F�Gw����*O���S慛��D�U
g%:�'N�8�7��b� �@��������'r� �Tϟ�D��86�\z},���'��H@Sl�{2 -[�EP	w0<�	���ɕ;�)
5B��)��l�1��B�I�D.���s�ۜnf�ica'�m�dB�	 w��s)TN��)S�$C��>
�T�S��9` �����ّK�C�-@���%A�)�v��fӃ*j!� kG��ɴ倍mD:@�H q��s��tS���&��4�wD�U4��b)�O����8@`��L���W�p���P�,I�L$,�N���Gؼq��\�ȓ=�\8����<���3U�9r���e���B-�=)<��㳬�>{d��>��$ <O�p�S��z]3�A�T�L�"�O��TR�n����%�
Ȩ o~�<���4}��kw�B��s�.WE~��d���(�� �(�)K�]W���.�1,�����'	��',`�	o��h!g-H�
��)�O>��鉣��1�� ��/��$k�Ȁ�K��,�(�����ڑN]�F���p��W؞T:���?\2,��2��L���y1$�8���V-^(a��eݢ;Q�8�*��?�.O>��Ĕ
H��<���v������ax��'��O�+���Z�0� �	lp� ����wH<aqM�W$ZS�
L$A3��J�'MaxR�..@��y��8S����y����od�!��o�8��Ν��y�]&W"ƀ�6@Q�l�l)��X'�y���:Po��&F�=/��Yy`�4�y��� I�����)l�8����'
ўb>��1��>\�U����6F(��꧉0D��X@Q,2y��9@�N�T�h��.-D�`듀I�'JZ�h���RS�YE#*�O�	-Ic� ���%� � ���hB��3�t#�Ies��/у���9�I� %�B֦��<{�@l�C�	4ȸ0�B*��� WH�,�b�,�	^���ae�ѻBj�1.��!RE���p�ȓv�MW�g�2�1��R�d�� PRH<����$a��L`��S�%N����C��8�'��	k�։���$A8Ap�kF/Y�&B�'o:|H7���%+U QFF�v!�C�ɋ��Ш"��E�Tx��6B��C�I7'i��"�ȁ�!l�=�'�UGtC䉕s�t
R��V.�-qs�R��VC�ɿ<�	h�#��J�`)���I�"�.��6� *3��m�ыذ@<�C��5L�p(:���4�µS�i�*J�C�	0@)�\2��9{�L=)`d�(<�B�f�v�SA��*F�tB�(T6��B�IkUTdj���?\��'*�%����?����Iv�*��/NtH٘R^!�ԤF���C&�� � `�ԥĊ)C!��
�nc�nPX���
�!;)!�³h?�H��ʸ��L��f��Q���� �ҵ��mV�'0`#�H�T�JC�g��I��&�2�|��H=0'���0?��M
2L�N���σ�N�p$��@�'��?�Ɗ�$��Uڱ��RϦQx�	;D�4��N],Ke�)�����O�^ā�n:D��skЇ!��]�f�@� ��N,D��椒 R�(���7l��s�)D� yR��e:n�bg&�!GY�=���'��{���'B��ʇ
�HX �X ���	���$��D{��4�W�u
G��/�#���/�yrK�B�u� l�C�C,�6�yr�y�t}*��A�N<�9���	��O �~� oEL:�t`�M�"SPMXf�ːM�!�$�?CfH�v'S�&�}Sf�7#�!�	�'���7�F��Qp����!�W1�� ���� �gYt��'ўb?M� ��'��!猖,���%*=��ȟ*��$�!S���EM�/o��`"O�<�B �r P��p�L��s"O�s�_.�t��sΈ�c���P"Oz��6&��8��q�D��	ӰiTў�R�'��	 �a��sT�L@$`1�f���'f�a�#�f����	��PZ�O���D�&(a$�E*Q�8YZP�$,���PD�t�L����j`�ͧl֜�P&���y
� f� �+L=ZX��e©@׼�0T��*�S�',��ɰ@� -����o��I�&��ȓB��,�8 �F���@��Fx�'$�8w@ۂF/�4O�3!�k�'���Z�ˁ5/��J#��_�v� #n#$���Oƿ}�F�3�O�;�D�&N(<O��nZK̓��pXa���x ��d-�(xBH�?���$t��3Ė�1!�� ��M�=���)���� dPbٕOz�H4lO�O�!�$�(Y� �Kd�'gv��jf�[3L�!�ą�@�:�!V5fh���V]�!�<C:1YT�ֹN�p���3!�D�"b$��B ��4 ��{��2�!�d�%��I1��_�=�bŹ_���Px��y� ��2)�1�R� �L.���뺟܇���P��v�J��� �N�/Ϙ��Db��$� ��K$w@�(�Û*h3�-��+7D�L�G�d�d� �M�$i�Q+��6D���U���IOy�2�u'ji˲�0D�|r�-�Q�މk�a͆^gd���+9�IO���'.�2Ȼ��L��>��I�3l���n�V(<���>kQk�1%t ��"��P�<y��_�;������fJҜ��I�P�<c��9a\8�(������z��R̦M�>������d٥_1��P�0@?&@�q)�a$!��ƅ,�Z�ң�J�5,���P�8��I�O+���F�Ō7/�� �r?,C�I��P<����,Ol�{�oM'��C�	�N<�!r��f�Zd�EoF�(n�C�I]Ȃ �Gڂr�6�;��*T(C�I)uR��`���O@������U�C�;��\�%��K�<�і�ՌT�!�!=���Ȑ'�+C�oda��)b����ᄘ;d�Yҫ�y*��ȓ^�DȄł{���*s��!�>=�ȓ'�4���7a�b�B�蔲L���ȓlW&�b��("b��p��Ńz|P��dD�X�6�ذX�Z�w'�(1ʜ,Γ�hO?�9c冃n���XR�I	�8���$D�P���`+�2a�;_�8�Bj#?I�J�)I�Z1-]��pA��}��Gy��|j�d��Lk�ĕ8=���u�_�<���]�Fֱ[��F1l��И�^�'�ayBD�3@R���T'X.���9�y"�!#��b	\rbA3Q�$q�\x6�;�S�O�NŰT��
On�B��a\TRד_���	N}r��o?�x�oنD;R�e"K��y�#� _�^p��R65�i2�B���'�ў��Hb�E�:^�6q�U��(�&-�"O��hSFɤCH�8���A�Bt�� �|b�)�(o�xЈR�?�L=��ٿ2 �C䉱�h@,ǚ5����SoY�S_���~��'�̹���A�R}��M�V;����u5
(ZS�D�E6:��F L�<���'�d|B���(b���c�y��y����O2ʓ��S��*i1��O��x�EFI�r��B�	%��yB犗
��ě`Z�VWʢ<�˓-}�q@��3>07f��H�� �ȓ�4�(0�^�xAJ� ��ZO�I��2Nd�g� `��m��\�,��4f&�J$M#PҘUP�m:�ꐇ�T=��*�^�2H���q�ǡA�����~����۹s18�SF×Gv͇�=��A�S�L>~^�Y��)O>�܇�S�? �ʂ���86���fM�Y0lm[D"O<<p�d�>���Hu���"O
������;L�Ձ�b܊g��UІ"O>�	�BP5k"��Q�Y�x��f"O^��A� ۀ�sAk^N��騧"O��t�ۂ+�p�Ʃ͈���д"O�t�`�y����G�	W�82�"O����#Ŝn�����7N
AXS"O��K���* 7�#Cl�4p��S"O�as�Ď�5�D}CRő0�}�"OH�A��
_���Wx/̠ �"O�,�G#g��g��f.(���"O�تeF��]���IɔrN�qU"O�T�w�W$�г�\:4�J,� "O���ރS��9R�L��Q�5ha"O
�� �ɀc�`a�T,τC$��R�"O�i�R�\�Xe�؄���"O
x'P����-n�����"O��Ȟ<+o���wPDJ�"O��sv��0qT
�i��l�����"O�"0��V-#����"O�e�@+���<颧B�g�6�˶"O̥���"zŚ�����.mxs"O���c�>Z�ĳw�])q�)�"O�ZC��M��y�.>Y.9�'A����̂c�8�f�wɦ�����8�0=�ȓ(Qp)Rkߪlo���ɋ%�t$�ȓ�v���iR?|~�Q��j�R,�ȓd�mq��"��!�(V���ȓ{�>A��B8ļi1�%�g�L ��I�F��%e���D� (�ćȓxި�{q!�:S��r7S�)��(�ȓU��E�w��&Q}�!ŭz>�\�ȓ�U���[R<�Qw����F��ȓgd�PK�W�@|�t
ѬI^Ё�ȓ0�I`�/UT��%*B�.*D�m��(�� �Y"�̔a�jQ&?{<l��j��=�h���fȫf�ȟ^�Nl���:l��ʚ�Nl�dĂ��\ ��r��Л,3tAR��N�.$�Ą�^�t������QV��JQ��Y]0S�AP�	(P)��d#��A��m�.��U�z98���h��`״�ȓ�(��O�(@����K����A|��q˒6�&�C�C�X�J���y� ��HA�H:ƽ�$�\�q��Շ�~��@�E� 7vL�V�6~,�ȓkx�����[��U4b�)6M�(�ȓ"M��А%�(�V��I�� ��u��t�!y�j#R@cR�|%�ْ"O<���&�������g��D:���"O �r�A^���"�L��Js|� @"O\4s1M��+赪��v�Qj%"Ob�+`��=p��ppn�>#�"O�����*k��U�p0�╚�"OVQsIH�K�FU��-]�C|,�g"O!s��'O��Ik��nc�[T"O|�#d�x60�ŉ�̈́��u"OD�0r#�=�h�ڡ�͔�*-8�"O�y���Y6l|։�s� v�ز�"O@�{��
ĦY��ǎv�p1"Ot cMڠ�jQ��揥S��lJD"OhT���Æ'�h��ѼK�� 2T�D���N�S�O!�H��� ��"6 U��	��� �`h%�h��̡���C�\(�xb���#����	4N�X-�Bہ>P8U�C ����$[m�t����N��Ɂ!�řj�i���xr�T+R/v�Hʃ-Z�򑱒���OR�"Aㆳ��O��u��꛹J��q�$a��$�F���'�A���&O��"	����O`,)b�����H�T.A���	V�#L��󇌒M�!�$�-��t�{&x)"�($.��'�F�j4f�Vx��ؒlܤ+���q ���T��J�.�O����,F^���L
��T&N6~�.C�
sN��v�R�R�����*�%+P2C�I*}4���iJ4�ڽ�LKl\,B�	""6q�G����rvc���C䉒z�.�YpO�d�`ѶIKv��B�	�h��y��nMo��|�%�	�*~B�0A�VXp��R�-Mp�r���>'^�B�I�4"�
@/_+�8�� �1�h�QsA�h<��*�U�z���������VX��b�kٝj%�'
��VA�0|)�����!=�� x
�'ZL��!P$}t�yv���Db�81I<�R��%x���b?�3��n���������LY�@,D��@B81頭@tE��q��0�vH�`ܓVl|c���x��	#��HQtf%��!�g����xR"H6W<AdŝkOP��T]$z�L��% S��1���f���@$�Ǡ$s��s.+,Ot��������LP!��b��I�*ҷt��e�ȓG�Vؠw/_��t!(����q�n$%�(0��n�Sܧ}��X ��A���R_6-���� {�lB#*\<0ǈт?Q���ȓ]�f)Q�@�' ��1�>1�&4�����l��6~�'��&!�n��ȓt�\�[��G>jc��3D�!7��j�5�ɵ�H����(�|Y�Î�?PΐC�m�8
%C�	+�~|��ǘ���-�R��)ei�A��Zx�7��dP�Q3�{�����q�0|i%#�\��lH��Q �p=Q�A!8��U�Xp��ɁKCv4�`�/er��B�| ۮgw���}&�\���T*(�Wa�`4�1�B5�I1��4B��I �6�Z�� �S�7	̵2�h%l`0HJ�=����
��p+�D(
�#`���F��Q?p��K)v�k��xܓ��0Q��6�<��!c.}=�����S�
H�="�H����R�yZWNm�<1bm�ȍ(�;?��`CCn��M�4s'�(�`N=2�ބB̈'�u�9O�8����1_摘�d��p�xak��'��܋3�>��xe��wL,6�M�g嗭�}��߭t����2C\|Yf��g�'�����@�JA(��P'������;��ȗe��J��(�C*čw 4�1��N 1�ݰ�)*;�Z�@W 3�O|�����I~���p�e�ΟW���у��7�IP"H�S�J��~2w�ڸ� B˹z;:q2bd�b�{9>y"r�'*D���������sT��O�Q҃�T+dBhѫ�<Dt���Q%�H�*�qq�U^UX�����85�����oh�}�u�5�8�" с�X�G%4q�6
N��M+��$��d�f��A�}x2 �*΍xF}B�c�m���Q:$��
3 ���a�>�O�	��o،@�<u
��D7�Z��cj�5��i�o��6�H|s���?>��Q�ߘ��S�OY�]	C���<��l`&�W=�� ��D�`\�I)c�&ҧn�� q���v���C�H
��q�Oh1)6��
x��Y�r��lG3:N�%�`� /@^,�E�/(�x,�ä;}��I�
F��ٲUn�<bHt�W)��_��e�P�5�H�#	�'���sI^�^��5_c	�'��}��3%�fX�'�����o�R"�!�O���ґ#�	B��ߢ?ZPk���0>�b�"����'�H�6w�}b��� 2�"��Bݒr�����69fbCjC//�%����>-��3�p
�@U>ɌD8v!	�`	8d���e1"�|b��h�Π��Y#6t�Y���y�$�3D>b�Rӂ���0<!�j�O�)��N�3�p�ŃX6S�x�+0D�	�ҧH��m��G�ψ�аA�8O�6Ԁ���4'Bj�8Ь8��+�e�{Lj�Uk_f�b�H�����U�&ѕ��h��x�qO��   �‣LJ�y�*��g�X	���'@�)����H��]8H���q�DU�eGx�|�h�K�J���SE�>��	n�zIe�a������C�'��!��F	
o�p]#D%�AⓓR���c��	&8|�W�X�3���7�(}�D02b�9R��'���ǂ �B�"<�g���]�F�I�4<�\�q(�d�B���˼���r��'6����s�υ���3���<��iUg[�:1�D�1.-�O��Q�a5r��tN��Z`��t�,}�i/[��p[Chf�!�Ѕ�;��i:�>�;fQ`��	�e(j�G(&���A�':b,�B��������1��vppp��,91��� �MP�O�>�:fohԸrr*�
oc:�p�I%�z��h�6MPdP�$����ܐ�	êV/��U�0�@9QiH�'�`钐�^� �G���TU�d���M�W3&4�fƋ��d�g���A�5��$ͦ>(��c#£�uǠ^�z@J�`�lF^)�qk��Я"�@����Xs�lܔ'��{b�D�u*�������פԩ.T���7*���u��!�Dm�b�R�9Z�#[�Xt�;�*T��j���)(h2���5�Z�!�W؟��Q�Svv��a��x����W�ةCX AG�9+R�W͜~����p$E�vqz����b�3Fl���T?t6��CΧ�|P����Z�џ���oˏ;�@�'���ʰG�/�v��(܃/�YaA��T�&���0-��)��d�kH"?Y����u�����U$P,'��!S�O��#p�ȠYL:����N9�����?e�A������%O�<�N8��銱PQ,�`�'�)���*�`��ȰD�Ԅ��g�O��� �R��,;��̈(z�9�O��T$X#koH\�;?�`R��yv�e�P��uu����?}�x����=D���%�#�<��q� �d��1�]P�(a̒����f\�F��ٝ'ǉ'!`�;ł�x¢��cn�$uv!���H�C��po 9�����8�b�ѭE��&aZ(�q@����`�Hxl�4_��@b�ڳk�Y�ek��M���fҘ�FKW�`��	�f�@xx��� m�x�n�#2��$fκX���W��%M�V��%�?�ݴ�p?ٕ.�?hl��"{r��U�^�F����b�§ �YьQmZ�3�iM�D��0�K3�y�#T�Z���G�`��Y�B$���x2CH"QHM��"̒j���7�t7X�A`T�Mkb-x�K!nǃl<���$�����1�v8��'�/~H��X��x����a@��c��F�"���#�݇�
P@�,�_�*�x� �v�V<��/�&K����*�B�HA����M��Dɶ�R�>��V���s�3u�r0��ːw~���e�v�P��!o��к��rs�P9�V�E]t�v����ǈV5`�:���",� �L�)}���&,�Ox�$h�x�7@��8f�h�џH��+W9r6�Ƀ�%?#r��O�z�ϧ9b�|�S2�fq�d3,}#��`[Ă!O�9���,�2@��+�tǎ11Ʈ*%��lC�+��c',�g䚀"� ��ܴs��'vh����U<1�H(P�-&�{ד�	8r`��F��1F�h�*֌\�1p��R� �Fr�[DIF�`�����0=�kRB |s��T-1�q�s!�E̓1��LP�"�94@��U+F�:S��7;��St�Ԩ��
��J�Ģ���9�'���A.@AZ�IǗ�_/�觡n.�"4�EUutYХb��>�r�ϿCJ�L����I!d(��D+�gh<��F��HN6�읳�E!0&�Qp���$%���šiZ S�݅�F|B�	d���9�/
)c�\Bd�� ��<1�'�D��B"|�H&�Z!zC��>te���/)㪱���0�O�8�%���,�θ�5
V�(gf�q�I,\$� ��[,�y���M�u�8��O]
܀Tk~!��T;5`��N" ����� Ƥ�y�� @��0� x}��9Or�
��H2B���˵OZ6"����"OZ���k�b֪��2��%���Q�2O���-�)�p�@
דdH�!bTaW%�1̍%}JD���Ɏch<��B�3&��v�T�>���g�A���㐊"D��cEmʰ٨��U�=�<�+6�%p�̥0�jZ�
$��|�c�4\lf���ǝ@����%�B�<���LT�ěv	@����8I��Q��J�h�ɧ��R��}f�m��р����g�6�y�Z$?L�����.i�$ia������?glt�@C	3��<���Ĳ)�2���{\���QM(<YfB٘]�,�+t���L��GAG*NB�-Op���l]�5�\���-bf����(O�83�FM5�� Jqj��D�Լ	�"O4br��,9�ҺU����P�8b��)�'t�
�����%&��x����u^5��S�? ���w&��u[Pa(���<�P}� �xBF�a��X�[�+����=	�Z1W,D����.ʚJ8X"2�óZn=pq�+D��ӱ�]:k�ؼ���>R^|�9�o<D�x��!�3�f!끲2PZ���/6D��C��	�s�>y)�4!TJ9�!�1D���F��=R��)�:D�(Az(D�8b�G�;I#����N�%�}�4"D��󑈐�V��a��d�&dXƈ��-"D��age^�G�̬���ȮA� !�#D����.�hE8i��fӖ{i�\�T,D�Cb��,7���53��8���-D����K `J��4�ÓkfpI�(D���`z�H����a\ #�2D�8q�'Wfl���A���&���-D��q��7$�I���� [F^��& 5D�2Saʵ�Qd/�!@R��`�3D�x˨L��)�$���m�>�;#E.D�4(���5 v��q$÷j�
�!�� D�,x�
>L�������<msM=D���pD�/e���;@/E�T���+?D�ʧFASԐQ�Sc$&8�x�7I=D��[]�O	�aĔ
6�0�4�;D�kc�%���`�fY��xQ��%D�x���ZR�"I��nL����<D�h03�E���p����J%@q�`;D����Lǅ%�P����#+| ��4D��y�)]�`���Ŏ�J2̣�B2D�x�!̮>C��7��"q���V�3D����H�!!`xf��0H��u���;D��d ])0~MJ��#��ƍ8D������~Z���"y#nMC�l7D����&n�6 ���+�^9��;D�(���=
$�<�F��^1UR��%D�� ���3�n��m�<%X!��"4D���䅞8�� �g�@ 
��DK`@3D�0���-P�Nɢ�F]�@	����%D� 8��*Vd\E��(NB�Q��%D�h�C���\�cq��B��� ը&D�:/�/ *E��H����9��$D�������>�j�� {���3ҏ"D�؉��e�f��'N�M.Ԩ�ĭ D���sʀO��PQ$ Jn���e� D�|P�#�o:P b�%!)���	��,D�l��*6��:B��B-��)�-D���u�S�"'�����=v^�Ӣ+D��S�O֚n�l�ѥ�/)���+:D�D�׬�*W�F�"���W��6D��1��b���F0S�<��tI#D���Wh��7�8iK�?C��+�/>D�ܳrMb��B��j�a#�`9D�< #)�e����%�Ԛ}� �b� 5D�,Iv�,���R�c74���5D�S�"�(@�!&��HS�be5D�hHwC�,O<�pQ�&%� �3D��Ϟ @�^�JP�ݝZ���)CG0D��y��F6_��A�b�ݪ+QRв)-D�h�`�K	�9UCF�c�p�T?D� �g6;�Q�[�dP)�e�+D���hR=]��(�
��}��
'D�r�(ȓs	��;e	��W�5z2�%D��2�
ļ7�* ���gA@��6�&D����[afQ��A���s0D�����H�̈F-�,Io/D�� tYA�eʿu��������*"ؒ�"O4�3��N(q��H�$Aٛ�x��6"O����9���Hy؉��"O��5��xБ:�J3<��)��"O�9C��ۛ'��<�.�)�B��#"Ox��U/�6��	J'��!�Q*�"O��R� �.P��0F��s���"Ov5��L�.��%[�$^+%	�Q��"O����@�)����#UD�R"O>51�'�(�1�,ڜC���#"O�(�,��o��d��MOW�n,
�"O��{�b\v`���6Ųej"O�$Ӷ@ܺ�\RV*ѱ"� ��r"O��tث_�`]ڢ�	8�8*F"O���;2�8�ѧ��VD��d"O �0o!,���@ϵGM �ٵ"OV!�@�݈p�@�C��W�
4у"O ��l�-!�=���Cg�)��"O�����G"T��6����Z�"O���b�$|��q�C��g�ı��"O�l���]�0�UHQ��xิ"OX�)�EC
m"���G��t|"�9�"O��`���v����R�ieF�"O���Vj�g��BC ݭ2H��t"ON�"qƈ�h���os?��Q"O�|p���'����`NL��� �"Or��c���h�f�
F���>�� rw"O$�TI0!�tq���RrJu)U"O6t���]�&���t�p�y%"O�D��E4)�z@+���P�MyC"OT)X�jՈM1���$G�]	e"OƭQ��-&ɂ��2c{>����"O(#�� +�������tBPX0"O�]�ď�D�p��C"Ϡs\��2"O�� QI�8�^�� ��16.�s�"O��1aK�X�5�w%��[h��S"O�E27+_�JNΝ�E�C'�D��';��p�Ö<o`�wo�����H<ɢ�^>b+�b?a��š�^\���?�d�GB:D�@"�A�DuS��ܧCoH9��!���Cm@-Ё�,�3��Ȋ-�4�+&��~�ݰ�iY�zka}r�S�_��I�E�9(;���,xa��O�a� ũe��+<����'(����T%@��u�ҤB	T�Zp��� 5-��9�g�$D��]��$�I�IŢ1MF�X�O\6u(
D[�
�)\!��m��U1�� �vp��J�<"J�x�J 4Q��4L���3��s��Ԭ8bk<�!\�c�L�x@8D�pi���6U�¥+"����B�d+aCAч.V��
2N̟(-��3�k���toƙډ)`*ژ�8��ɁQ�҄�iI��n�s��=+¨����=�D�A&��7��ś�'V�qF�Ɩ7���
/�B0���e���Cl��.g h�%?����{�(���(����Q��K=G���O�Y��˽ǰ<��+���xsԭ 2n��az��ҹ^�L�wh�D� 8�fO�'E�.�G�t��.\$�y�茤�lI1w�ـ\���bCI�V�����E�
y����?Q�Jh �ǛZ�l�!Vn5��J���l;�=����x�vӧ���G��b�+�
J��eH������$-E<AP�@�u�b���@SUp� I��9P�\bGn�6Mpeg��Q��I�#�>E�hB�*��՚ק����'(^��(O�}�G��(��#}���H�Z��yh�$� �r�>�D�+:E�)�A�2O�P�� �k�tkKV�MRh���銅]l�F�W1��)ʧ5�0q��(J Ј�,B�P�h�!��)¨��@"���Go�)jq��%?*�CH`�h@����q�S�ċG	�	���P�>�5 ^���QH�du^�hG���:=,����A�\��iZ.�"��-ȤO�0��Eh$���: �O"m�a�-G�,��M��}��[+.��L�#(��|�a!f�A�'"��`����S[6ME�� �T�͆Ҿ�`��צH����>���.N��-z#D-O쬘�懏�&б�$ţow�����*ff�(1�B��)�'x]丰���p0��P�4�h�"eF�L�a�'V0d@��!zr�dsf��6Od|2�'v��4c�2d�'�<��OO^�d�p�*��G0{HH�uN4Ƥ��
�Cr�YV-h�V��ؐ]�LhGW)T����`���	;;�N�����6�����5�l�7E�DL>�<I�dӒ�>���K�7�b>Qh��LM�m��S]��P �1���_��	p �1Ob�)�O?`}���32T�l`�i��!�'�ux�r֊�M?E�4`�9���P���f�B�zc0W�H����f̡KZ�J0qAΒmب��I��@��'РIy]w1�Hʅm�!���O�ٲ�B�37�Y5�5�,U��a�ҳ`5Lڤ��~׶͐�`���l��E̢H=���W�L���l�Y��	��T����&�M1 H�"pǒ#?Q�G�?c�.��,*�I!D)�	:���$Qvm;ń�W`�'K����j�"���Oi���(R�����*z��A0�Z������&B�W�>�|"���pD�ȀP�p�*d��;�x19G�@����K���6Xfi�h��'�Ԓ�OQ4"��	���O-��Ӻ[q��8����t��:2L@��cy؟(3�"֜7of%jFD.ȶ0�͙�`��!���gU@��Ҭˢ}ܐMv�>E�F�W���p䇖f}���B����O�U��バX�c>iC�W�r�����m���`�&�䗉o���@�'&O�xA�
��@Q���TI�2@ى"��\y3�":`�&�b>I��i$�U��`�=Y��HsJ��'u���V
OV�S#��G�e���j�Hm&$�x�I�k�By+f��|"b��5��qb��
X�:�aF)�x2"ؕ6�|��]�Cl�Ыѭg�l��+,>ޡ���5Hr�Mbw��� D�A��&֑u���$�`D�,q"�R���Y���n$���g�
��B�	�)�NA#eS#w����9 �v�C�t�3o��qE8ӧ�|����9�f��B	�L�����"O�t86K�+&��xڳ�=�D��R���I�
}P���1�3扨S�NX�*O�v��[#+�ODB�	(Q�ZP��J�+_=��{�E�c^R��'d\������'OPx ի�/n�*4zc�˵���3
Ó_apQ����HY��'Jb1�Wj�ih�l��޸m��P�'�$�)@& TFf�ad�ٹ�	R�O���(�2p-�!L�"|��C�-2P�գ��m�Jx���H�<�&�Ŏh��EӔ��	=���w�o��'���'D�g�<=�|�f�� � g�
\`B�.G�D[��G�.ܰ�J�V�hN@��Qȴ��b�@�"�4P�7��2yh�!y��[��y�؟x>�T��B�xʺ�Q&Kɗ�y��	�Yb���O8~1r���W��HO�}�����h�����I%�*���!��1����"O>�Q1!E:X�hH�M^�v����2�SX��%��F�)��Da�j �i�xM�Ɯ�h�Z��V�#D�����Z�c�$���+��w�.T�V�m� )���z��Mi��'�١��۾F�"�ᶋ�'(*Bz�\�2a��љ�������
x�f+��$�� R�<�GU�l�u�C!D0�ع���d�'[�e҄����G�����QN���;ŬY#�y2�C�>�(��祌�J�,���"�'�4h��mS�}Y�`�O?��&N����CZ�4(��A.J�| TB�I����T M�~���ɂ(�5L�I��7LL.��zB��/Ow"��p6n�tO�!�0>�1�Ƣ~`�����j��a�g^��n�Vl�G7���ȓ}/q��nN�Q^�����J�B��Gx�5}�P(�r�\�O1�ѓ׊�7:�=����;"R��p�'n͠���!G��iЧ���!��x�f�Vh,�RDo8���O���Ō4ܭ� \DQ�ᱳ"O|�2	Y�w/X$�t�ҩSX8ŒF^��k�bѧ��{r�xF���"0p8�p��愼�y��ԓ$�4�H��oа����y
� �%)'�ٿf>
��鐿ir���W"Oj���M ���*y,	�d"O�D��7}�*�:$|��"O�<���d���;�&�6i�0ۤ"OV,�T�� !�6-1�e��L\��R"O�1#A/�"���TD�"z2��"O(,A&�M$LU.5"���!?��"�"Op4���]I s�$ ���b"O�R���*WKh٩�J�9�D��"O����,��H�)��)QU1� "O���h����(�����"O�0U`M�!�z���X<�ܱ�E"Ox��WeU�H�	��fMj�(��"Of]�W��"Z���1��RD�:�+"O�l�����x8Sd��/�`U��"O�����Ϛ'+L���C��B:(�"O@�a��� x"tj��ʰ"O��;W��g��%FaZ�_�0�[�"O(��)B8.r2�z�������V"O���^7^�$����K1h{���P"O`�) ��5]�<Ҕ��.B�+�"O�����;cn��I�;kl1��"O�(�A�"���q�ѿ
_@ٺ�"O�����i,��w ԙ0�d��"Ot�Ӥ�P��� ����:�I6"O��R�.'=��	d.�+B�1�V"OZX3��N�.�:���L�	�"OJA���)��M�X �T�$"O���aLS~��!�J�;Y���"O81)�
�9�z�f���Bb"O�Q%�V7d�6�q��c��(X�"O��Uj"&�R�䲌�C"O��/tr��ր�*JHa9�.�9$��~���9y���A�A� �ִQa���(����N�<7Ĉ8]���c	�Z2�Q�MTu�<�fĉ
I�2�`J�2b�����q�<���G�(k���q�LL�tqU)R�<9�H�X���� h���(��MF�<i���'."��	a���;E8�G��J�<)�,��g5T�́�gK$P�GG�M�<�5���N���c�c�83�T��	�@�<Q�L%&��=+�K��H9��{�lQg�<���Ơ|��U
�+=@���CU�Hd�<�e�
j�U��MG�&.���֬�W�<��h��{'\D�Ř/�N�+dm�m�<A��5�F@ ���^����v�LN�{���r^w�,�P#�T�c��4�p�;�M�+Y����'i�xgnۚW��O>ux��Y�!J��PG��5�t�a�n�P�D؈u��\k��>E��5`��U�t��)���3�_ 6��T�/J�z��OQ>��6�:%�Aj]ˈ����<>�ɛB��dd٭O���o���0|C�]�$��8� aВ����QATy��AJ@�s��1Q�IS�Of��0H�~׀5 ��¾҄��AAb���g-�R9*���h�*��^H0��_n��l��F�J �1�!C�a����69Ol��O�0m��Oȃ*�R��S	�D�/�^��8��'�<���i����z� L�A���SĐ4fk����" ?9�ȡi�Ԉ�#C%}��Ʌ�
�Q�B��}l ���'\:	��Y)U���&P����|�=���׾�X����l>f5��i����`Uk�S�O�NƐ~�z%me< ��4���k�fq��>�$Q�K��B�6 �3@�gbiq"OnL��&�3l���
a̪	8L�i�"O�A�a�
"��E��0Y\��"O�Y��Fw��h �%��1�C"Ox+���?����N�S|�(�"O&��A�3�����R)�%ۦ"O� ��e$��p@��O H��"O<EspcK ߠ��r�ݙ �E��"O2I"����Zh8��% p�tM�"O�K�mZL�v� &#ܾ}�84��"O�th��[ ���X�� ��42'"O$��B�x��Run��0�J�"O~i+�`�$
�I�&��X!�w"O���'օ_W���kų�(��U"OI��@�8Q�:�*�K�z�p��E"OB�9"gԋ`.�5k�L�	~�TJ1"O ك�5um&�+�0Z�p�3"O�}��A�=m;"A��I�X��Y��"O�Hd�([�`,�)+V�*�k�"O�Lq�Ա1�Zu{�m��r�@�P"O@�a��Y� u�@A��*�X�#"O�ȧO.b��kU��?
м�e"OD$4`�m��@�?KҔ��"O̅@��[�G��@��D7Y<�Y&"OZX�S�[�)w�Q�1l։y.z�Sr"O�a���4u�l�y�ݕFȂ!1"Oڠ4/�~�^�k��@(�@�1A"O�J�L�ɸ��&]F�q"O8M��M½��РFɒ4W�pW"O0�C#�K A�2�"�×� =��c"O����-�/�=��l\�����A"O���g�0�@��),*�Ή)b"O8��MA
~$v���*M
**F܋�"ORyy�D�--׎4�	��>�1�"O�!���}���z�nױr��1`3"O`���W)9�l�H%�1�h�J"O��X�зb�
�"��J��!"O��bǑ�&���26��z	|��"OL�P���N�"�X� ��|c�"O�XhC	]ռ�yQ�Z �n$�v"Ob$���O�f�8Q$\m%��"O��ߦPWƕU�Z�Rd6��"O�]q���oR�]:!�Q!F^���"O<�h�B$ H��.�.���"O&�Be"@�躥OJX���Ӳ"O� ��p*�B�,ܶa��	�
��B�I�Qh�I����-��Ӗ�;t�C�I�o����pm��3��M:��_�!΂C�	@�$�1��F�ƀ�P  �VC�6)n�+�� '֝�Qφ�C䉅=�n08�H��+�aSlαr�.C�	�,���KD̑Q	��a
"C�IN��݃���(�� gDP�	U�B�ɆEM��@v�H nU�2 �&'�C䉊A�X(PJH��QZR��E�BC�	-(Q.x�u��8,K�"�iR(ID&C�	f�*��G*^��� �98�B�	&Uɼ�t$�<G8<]���*��C䉿F�|I�p X#�#��0,?�C��(@�R�b���)��_C�"B�I6Iՠ�S��N�&BU�'HZ�K[B䉙&��H�M�k�u�W���y9B䉼:��@0�bŽX*�Y�Q�C*��C�	�A�De�:t�a���kM
B�Q��p4%��H`�d:y�C䉫yu�5�J�h��Ԙd�>D[�C䉿J�QʣD�9e�� ��4�C��6e: zԅm>U&!�b��B�	�?��	F�͡R :ª�:ϼC��	r�����iE��	�ĝ�<1�B�)� x	��]`켊��=��M�b"O q�5ʂ�>��ѐ�g̾H~:�"O8R��Фs� �1U�֡;uBs�"O*��j�6�j��\�Kp:��"O��h/�:fȵ�5+�) q�<`v"O�A4L ��VX+�#�Ml^<��"O�Q�E�؜� h+c�^��J��"OZW�,,2�j�N6^(tSs�<�6+I�3�x��A0\�B	k��Qm�<��Ǎ%b � ����k y� M]s�<���$H���\xX
D��E�<����c��-y�'�	aX#*F�<�ÍZ<k>�$:���tOL}���L�<� H�s�D|x�dL�W\�,%!�$�9!��Y��ٍ/m��H�!(!��%-��`�a��	,Z�X��Jب�!�	y<a؅@�&sV����)�"�!�D��]�:���Ɣ�f&�]�g��	n!�ހ3�vĠ���?)������)^!��6���p󀐹u����:\>!�D�M݂T�P���$�^D���	:U!���~�(ŋB�$?�8��L	�!�ݩyn1H�f�D\�%���!򤉭_��H��S%!�YZ���7�!��ߍ�>��� �/(�m"P��(J�!�Ď�B�.�)6nӚ!D���0 
q�!�dxX��4oP�{1��D��7y!��,��h���i��5B�}f!���q������G}�:Y��ļ8�!������j��tʵJ&Y+!��z�8I�0M]�J�<ಒ`	�!�ē�/�����E�c�^=��<X�!�, � �a꟡Zd�q2��@2J�!��P��S���e���ۄH�!򄑜�xy���!s� ��� Iw$!�d�e�0�#��� ��0�`_�*!�D�����h"L��z�U����m!�D�%��5T��.:q��M��d!��{@�!�GI<lE�p�M�P�!�D�b&�IX���\f̐��H��!�$�>ٞ !���@���KF�!�d��|��EAԝ��	��(^�!�d�*$�Ұ�Ƅ<[D�`���Y&I!�d�)̪ C��o����:<!��K�N�"aJɅ&�CUoH� �!���y�b�!6镲�B9�"O
�^e!�F�܈�q'��Oy`��)T!�D��R`iQiU�[�<���*P!�dC(7tm��+��@=ְ�g�\ P�!�D�/�� �UN�Cj��얍�!�� ��z�l�a�"\��K���!�DO�K����Қo��)۷���
S!�dVX �C"-S�>�.���:I7!�D��+>�jG��h��4Q�_�9!�ز)����6�0��ѫ�C'�!��Aw� �#K]������8(!��X�V:,#խ�H���M	�!��V,.!G٦��1�=C!�$��Uu\�Z��Ɇ>�*4{�ǆ�(!��sϲ��Bi�f��}��B�B!��!w��DzeΒrv.��� ��H!��Đ>�\���B�n��	p��&!�!�dٞA
F�)6��Q	��X[!�Ę2o�,��I
�S�p�	7��nc!�� �`�AT�D��y�$��*�ڀ"Ot��&C�(a�Рѣ�/_���"O����#Q2bU��Zr`ڛ(fjt��"O�xkM�6$-ʵ
@@�
5'��`�"O�� g�(K��h�����Vx�y;�"O�$k΃w?J`�L�8Z�Ȋ�"On5d2��kS/kZ��S�"O~ɰ�gI�.	VMRu*^  ��dX�"O2�����) 
�y5�,G����"O���13+rt�c9Yእ�4"Ob��	َ8�"4kԃӯ\9��"O��*D�T�8(I�0��_{��s"Ol�0Q�_�^�@���>Ll�"O��%jݺY����'�́?4&��4"O���JX"0�� �̹�e"O���P.nv� ��l�P|�E"O�Y��������G�@���#"O�<�mȾuT�u�a��c���8�"O(Q�V��� G�$7��	�G"O�=yq'�:w7HMh��2p��7"Od`��+%9"������`�@"O��a��P��X(����2gT!��>,�#���#3��M{2!�ص'�})�fݳ_&��ْL�cB!�$=wv��)#�;9��p�@ !�d�-`�pb���9S˖I�4
X�n�!�$�(� <��E�.��5�7CS)'�!��~6nq4�3~^5�b'�!��)g��(���*H��š�v�!�D�d�ș2��֧0�h	Y��A	i%!��,����P#3� @*��߱$!���n3
A���:���KP��M!��I2kƥ���\3#���AJ	�!��X^��ꃀ��c��1��Z�=!�d�f����Xk~�\@%���1�!򄗽w�N��Ԅ��/�� ��7!�����9牝)f��p�� 2`�!��Ƃn7�T� ��I�Q�G#z�!�$D�D����b����A4O�!��<t��]y@�ɶq��4`ۋj�!�Dި`\=J�&�%^2��)�!��ˠ0R
��V��>A��0f%�b�!�+.��������ʄ�G�G�>m!�dS 41����f)s��4���ڠaT!��.X\���Ųah��#1��L!�!N>�PRb�)`Q(�C�-�J!�d[>a��'׵4i*4 ЂF�;B!�ė�@��I�����8�g �+!�ތH1�=��<>}���S��2y%!�D��ɸ��"Z�b��Ύ�@ !�dBk����fW�;~H�w���}!򄜃@�f4�eP1b�H#�}�!�A�X+�9�%�<��q�ve��$�!��׮8O������!����#�!��u�YQQ$#[<�{�舅:�!�d��/U�x���T�!1h;7@!�đ16b4�׋�k�4�%ǖ�+&!�$�.�,I'LX=_���W�X2!�D�{��ٸ'�k���&I���!��6�j `� ��z��F�^='�!�$Ք��䚆��h�͊�M�$ !�D�WI~ur5c~�.xz�%
�>�!���O$mj�H�"x
��H%�K��P�Sh�6Sqz)z�H��> `�A%Q�<���m� �'�	�Dȝ�p"#����,�OF`�  m��o�,.�D4�Fӳ��̉����zIz!��I詒B�'2*����m���Z`@n(�d�����?����䓮?����'���������9 N�f��`�p>�'u������)����7	ИB/�3S�+��,<�D�<�2��#?H�a��ߕ�0�˶q��̪��P��P�*}bAI-"^꓈?G�4F�}'?��Q��,Ɋ���a�4� ��(,O4��Ρ7�H�B��\eQ�(U�(�h��c�b-z�S�g���axRK���?��������@��#�Ă�NBC���O��d5�)��?^��	B ��TY~mh�L\!2�x�h���T?���kĽX��@c��� y�-�RH��XyR��Xx�a�'$�O��1�i,r$��D	'������T���G=ON��/t/�<-�1��O<F-Or<�[�m�r��PJF�l����x�X��P��ȟ��q��D��e�K���a7�x2��*�?1���'��'+8Lq���1��@	s��(_ЧO����O��O�c��y�f�e(�T @�8���'�k�'����n�D0��"~�u����#A8�
b'#v��)�b�`�'yL�b���i��O:=8��s��)�� �x	 ��KP� 6?O|��M0@�(��I�z�r�I����x�(�3D""�NI�TLɆM_F�+4�' �����0�3��P�f�� �W��Q���\���M��.���0�S�gyB�iK:D��@�7���q���$+��%�&��vX�����L�D?h�1�-\�z�q���O ̓,ɛց~�X�On������#p���bg��6�±�#��2}�;Be���@X�����m�F�O���J��`�R%B֩=!"eJ�E�o.�AiZ�aM����-T�3��n\.M�w���hJ�8'�Dh:`�Eb��E��%��P��
�r�,:2kݚV�*������p���M{����O�b��$%��?	v�E��_~e{Ǧ2}r���������Y^/f�Y�%ϯ�P0R0�|��M�`V6M�<����*Rf(����ߵ��?C�*��v�"F[z1�5�2�$ F�޼͓�?9���*<0O|�G�[�{�ʨ��C�R�ԲÊUX���6���#��1& �?���6�Q�]ky�ïP�&�P@%�< �C���˞A�"�'f�7mq�NH�a��N���JW�� �`�S��Vy��'"�O����g+��ߌ���lBi��`�&��c���i�6[#�e00�Qt2";��	^�z���O��O7md�<&���'�r�� ���   �  K  �  �   �.  N<  �I  yW  7e  s  �~  �  ��  ��  $�  e�  ��  ��  D�  ��  ��  L�  ��  O�  ��  �  ��  ��  ;  � � % � �  �& �/ : G@ H �P X S^ �d �j  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf"O�Ya��=!l���Ɔ�b�V��!"O�!)��Y�fx���eE\z0	J�"O>��pg�0Z�2=�C�A�Hy�"Ob\B��;h�`��Ɇ*���S"O�h�T�ÕZ(jܫ� ��+�Ƚa""O�A���I�{"��qReM.v�\�J"O�I��cR�G�Fm+De����(�"Ov�M�{�Ҵ�U���F�T��"O� ��M�g��l�a��8{�Y*7�'�ў"~rІ�$9�b�(p��:�� �t���yRI��Z��U`�� 1��)�#�چ�y��Ӷ=�
5 $��7&�\|��bӢ�y�/	�Km�s%�(}�E������y���\���9�)M��P	k��R��y"��9:*~��`
���r�:��J��yҨW%+z9) ���5(}ԀH��y���w��̙��E�zt9����=�y���g봁;��>Sb����y�/�$��e��E�|-�K���2��'lў�O<z���K�2v�����@�%1Zv�I�'k�끩Ĝ{y���6���,�|�H���5O
��&��2�z\{P�ם%\p�	1"OlU� [�i��a�#HB�br�͸@"O� $H����"�T ��Y( ���§"O�$vH5
kJj��UcL�ؐ"ONtb�b�!�&��"Ҟ�H�d�'�Q���M_�E���Ό�*C�?D���4BN�g$8d+�m�-	�����<я����X!Z�eWI�a�tHK�1:�B�ɵ.����C�1c��)��
��O���p<� �Q�?� `�E��Pt��u�\I�<��O3\;��K�&�mجU�2��~�<�diI?c��׋����!��r�'��FyʟP�i��V�i�䐰#,�FsH݃�"OXY��m�+����I=��v>ON�=E����M�~y�%/Bi�dgӕ�ybOAk�iξH2~ݲ4��yם�b�;�R>?����v��yB*G?A�=d�O AN�q�]��yB���t��EH'%�>��h��yS�R՜ ����Nj&f���yB�?ߎ���ş&q޵����+�HO��Ⱥr�y9�&��
 lHD��w!�$Z=��PE�%s�Y�G��]�!�dT�'��k6mY�3��Q$��)9�zr��Y�p���;0^����,[�!�L<"���j�oĵH��R ��JqOB�=%?e��$�,xQP0R�a��=D�(p� N����MІ1���跋8D��{���;��]�"�<%v��"�5D�|
��D�JF��rS�ߢ8�y�%&?D���ǚH��T`��.V�V�8�� D���DF8a�i4g]#"e8 ��=D�Ը�+۶}�.͂�A�e��]�t <D��HS �)������Rj����n?D���3�G�T�83������t*O��b���0��U:)A&p�ԁ�"O�l���؉i�*mK�j��
):�SU"O����CP^	�$k�L}&��"O�8��ԡHL{h�2~sp��1"O��s�͂����' �(g���7"O��0��[�`?j}FόBB����"O��+���j9��m�1b��xS"Oj���HқO^z�Z��<?Y�qJU"O,�I��W4�i�̀9Q�Z���"O�x�I(�f�8'
��~l�q"Op��/�9u�����e�dmq'"O�)RC��0F�A��è�qC�"OJ��4�ߥz�r���J�VR0��"OV�����E�!/c���5��Q�<�%Lȧzlb�.HZ�j#�O�<��ɞ^ ���f��A@օr@��w�<��I�'ub��è�O6&���r�<���Ӯ1hr	�!�έn�XM�s(q�<�NT&!�|��M��|⣀k�<�rS�ډi��˖���r�+�j�<�S;���إ�3r� ���p�<I6$��6p�jFD�+q�<�g�'L�e�cH�q�n�H�" m�<��j�$-j���c��%�I@7�g�<��`�P3�LB4�[�}�t�K�'��D�c�'ʢݳ��	ݒ�{�'�E�gV�i�L��	T�~d�	�'��I�U�Q|"L��b��spd��'s�!{��N�ޅ�L
^1�F.L��y2E^�a��(��(׸6���b��y�g$Fn��RL%6��Ar�ʌ��y
� A�W�V�:�=h�(��,��Hh"O���W�ΏCaN4g��	W$Is�"O�aa˯wV�� �# P�5ɴ"O
ygl�<o����nN�3�N�"O�E�����>S2���@�m0l�k��'�b�'R�'�2�']��':R�'���:Ю�t�z"bX̺1�'��'���'4r�'��'��'���ȷ��@A���nR+/ܢ�xc�'�"�'���'��'w��'���'� �!�T�YqR�a0�0��i��'���'�b�'���'g��'rR�'�(rDΈ����b�*�Z(�E�'���'[�'���'�b�'���'��Ԓc��Hq@��<��'�'���'_B�'��'"�'���'7�HMˎ��u�bJJ�[�n�b�'���'�2�'���'��'��'�䱵Q"s��Y�eb��p�Ҙk�'��'=B�'��'��'���'
F�k���$�T��Q�xI����'u��'yR�'��'�B�'��':tr��4��:vo�J.v���'	��'���'���'��'$2�'��S�����]S���Px���'�'r�'���'�r�'���'r��'|���l[��p�#O�t�v�'�b�'��'P"�'M�'���'醜2`�R��6��1PX�v�'|��'�r�' ��'�!$=b�'���y��2�HY#�`�9-X�ȫaH�O�h@��% ʓ��4�D��&�Ȣ��9�ZQ���A0P�t��'M�B���M��V���|��?y3��6l�'��1Ф�$J΂�?)��Ș\0XÃ�a�>X̓��/Z��Ò����	�BtR�p�!Ҵjl�Pq��#Z��j�P�0#I
B� �':��9o7��n��B閹"
t����|>����c�S�@c�H��"��5�w���aΐ�3j�H1jT)a6��%�'��Ǚ�E�B�$�Jh�ȟ��Je�!����C��E�Ѐ�&gm����9#A�Yϓ戕q���O<!:�c�Gy�9O&D��Ĉ/����!2x��E\oO�!���E��<!N>a��U����<A�~O���6�_�d>�� d���?I�Mc~Ү�>I��?����v�K�q�"љ�O� Qp�!�	��ml��%���<!зi��Ya���A���)�1�w�'6����H�L}1rY�%���NةDse�'��l��^���'���.xV&��r�Ҋ�P]Y�S�6E~�3)��b�"?���i�R����OD������j�xa
��	Jܜ�A��$�4e���'�0��3�K�Z�nY�i"�	�z������֦A�~�:�P1̓�h��@��Q�L�R�Ī<���'w����ʐ="r�'/"�O���h�!b�q0�F�v���;���^l�8<�d��b�矤�	ڟD��I�ft�'�(����݂a�t s���5@�|�Z�>	�i��6M^� ����g^�i˟r,;'j��J��ikA̜a��)��%Ô~��x:�!�5W���Qf�?]RT���o�5�`yy�e�O��ʱjͪ1��l	=z�0����즠�`�O,���O�d�O��:���(p�҂�?iF�@�H�L��@�F�t|1zU����l<�M���3;L��'���0���}Ӝٲ6*�L�`��!��[��֡ƣ?��-
�	�=�1��db,�ת��媟���$J����eӂ%#�DX�1���SB��D�jh��L�"�(p����?����C����{��� 3d�QҲ`�;fp9�#,K��?!��?�g�N�2��<ͧ�?��i����7�y�c$o;z�R틨m�����C92 9�'(��� 	�]|��O�F��A���p&%y��D��9v��Wl�  	i !�R ݀�1O6��7�j��)!�O͟�9���Ŝ��I՟4�I� �
-��7WR�h���=|J�H����'�h�k���Q���'R�O	��i��F�x �4#G�y{�IR����$�O}��m���l��%%��Ɍ-����46���O�'�\\���SR|��+k���鷍aӬD��cj���%���3���YӚ�iށ�:�čZ��i(E��	W֟���&hAV��̟�����xy�ս8$hUJ�K�2g9ؼZ��ڃG+��bB�Щ���'n�7��OR�����O�oڿ2�x�@'��:��p�y��� �4�z`����Ml������<�'�82~�}�0EH��c�lY�-L�,��b�Yr�l��%��<M�	����%
X����I��|��Y�(�O�(����9�F���G�1CZ"X2�+�x��'|b�'��4(�/����'746=��4�p`�>�2� ��r�@P�㦍�ߴM2���e ��.2�iB�u�A�>��3��(~1�y��I��"��U��7O=��,]�y�/��L��đ\1��d��@)����O���GCS���J!�� 7�\1�`�O@�d�Oz���<�@��:m�����?9��6�4���*l;<���J�,�D�C�ZV���'5��W��EgӺ�Z��O�JF�P�H ��z�(���p�M�)Wn�+�'.b܁�����foI3v��$E������'���� ��>Ś�o<!z��r�n���d�O����V�:��/�	�OH���On�B��Z�K���+0r�6�v��\	%��ɖ��O�D�香�ɶ"���Ӽk3���6�B����P�D�6���C�DD��6��h&�C���,)Bd~�D@#��$��ikp�$L�/h���`Q�r����iI�>a�\�m���b�1`�O��d�O��	G��;׀�l�j4��ϒs�~Р�	�<!��{���)O���� (� <���Ē�V�A�e�4z���D��
��u�'�B�i7���'ډC��Td�����xb�������Y�ch8,x��i�e�"=OT��c��y��	? ��Վ`�����;`�i��X<\c�����\�&}x���Q��D�O����O�Ŀ<y�E��j�H��iq8�"U�äGm:%`��:ԃ��b>���'z,@@�OP��'�.6MŦI�[3�����A��|a�c�̀7�H���\�J��$"�.�y�K��q��խ��y+��<�UB�ѿ� ��X�D0�*�8��\��j��+x�	�AA�O����O��I�!9����N��x��J�;-�	�a�Ͽb����O��$�/�θ��<���@����I�i�:�	�i��I9���8M��e�q�U�w����c���b!R��oz>�w��ssiM�8i�A�CNF�x�h���H(jpT�U�U݌����|��#������?��#�(�K���?��[p�3#���#�✚�Ց
� ����?a+OH
��Z��ʓ�?���ah.D*�#1˦�3����w�
h�I����Yʦ���40�b���\�&ĀT�p>�#�3��2���;)*!A1CI�vaRH�P��!C�,�Dr�� ��`���!yָ�i�iR�n�@����Sm�8V�T$���A���9!�.0�A�	ȟ�ԟ��	~y��P�VJ�Dj���z�t���DY�N$�FO5~��',�7��Op��ԛ�Q�O�oZ��*R�"<yz%�
�=Т\YشtF�q�C �>q��$��푈�?1�J7Oy�֝=$�1��<Od���k�%D��rC�D�2"ܨ9D�W�]@��K�&�HH��L�O*�D�O��	ǀ��ʧxƖ�CvǗ5W�*`j�HQ.S����H��Y �c���?Q����m�|R��e���wC+X"<�Ը��ܫ�&���T�ӛ��z�B�v�O��Ku����	�F���ݺcA������&tH�X5(Ϊa�z�!F�<�6]����֥���'����hv4Q��O��?1@DY�R: ����SG����JD��?����?�����$�[&V�c��O��d�O�Aa�i�>=� �)��OH����O���Ĝ�H�O��nڃ�M���W?���8Y�X�#�� k��xEA�oln|y(u� @PD_8"�fX�fƆ�!�p�	�k
�+�'l��BM;y�ܬZw*��⩑SOF����I������q^e��'�q�۟����L����	_a¼�ʅ {b蠈#c�ןP���B�UhH�Iʟ���4�?1`��{~�w�$a����(��8z%��\���b���MR��*n� 9��B�N��]):Z��A��@@�v�I�b��mWrU8��͎#X٘�E��5R'1O��82/�OYa���b�J��Oj�d��ұb�J�[�^����^�=��$@L���ʓcu���D��?����?���l����'�?	D��a��� eȭ
���;�2VK�Iԟ,nZ�.Z�I[T#��?e�ů �4zJ��� �T�9����f]H獢��	�^N�а�'z>-jS�n���� �̟<��ئ'�����j��T��w مD��ڧ��ƟP��؟����ܔ'S\u�����T��%°	.ZhP�	+{�p����I�3^��d���D^,j������O�6��T��R����C1���%�J(�v���Z|��`R�'�8���Ɉ׺����?�T�I/+u^=��'�"tp0�T�vQ�]p��5* �����<E� �	ϟ$���?ȓ#�o�sޭ;�C�0=:�3l�.�TAQ��W����	��䀠!G�|v(��ڟ$j�4�?!ŏ��<!�i�b޴�Cי��X{vRs�p���U�iYu���M�'��]w��fz��\�8jM8r'ʃ_; ��$ Ӽ1. R�j��?�%��?��ē!ETB���53V �酬�O����O���ҧW��]Z�#œ,FY#'/�O ���<��I7FP� ��?)������٧l*<(�b�H2h�lx@f���X��h�'�:듸?���,7���3Or(�'u>� G��T+�58�j��,l�vM�	O5t�(���Ϧ	�1�P�<�S&R�I.:��'��43���=�9��'��9+戉���O�t�Z�r����O���O���<���43�2!�ϕ V����U攇h�Z�A���%�?i�jn���'��X�Or��'C�`Y)(��}���W�Ee��8� ݭ'��*��MC���ee�.W�TE�'��D�ʺoZ�\͓���s�� 6�8�ك�ǔ4��	>�?�&�B=����?Y���J����)��ոK{�d��`��uh�
��!�0��O����O��)H����OYlz�-�3��>,��Qc�!�A������l�ɫ���i�����p�$�G�e��Q�
�>�*U텒	h>HYS@�rR5Z�{� ���4��1u�ʓK�gM-�2�c�'�x��p�L�(���G�
8Y�<�V�'\��'Ob]��Y�D�y�&5�'��F�m��%ckګ��b�O���	�Jc����	�X��
]�����Rٔ1��σ0(�d��b̪"
b��f�N���B(@��ӆ �j���6;O�ݵ.���7P&)�R䉯m ��yB�tl��?���?Q�!�/[��8�K~:��?���uҁ ��Z���SG���ni�Ip�D�}�6�^�?���7���'w��	�O�5��q3f�:�@�ddT�@��hp膘���!Cl<�p*k�e����<1�Oɐ[�ם�02��zbk���R���"56*AY���q��I��?�3��fgfP���?a���F�ղt���I<i�(�ǬƊ&��/O�i2tE�-4sZ���Ov�d��ܼ�2���d��C����pI�"�ꃰU�)�d'�>���?@o@?IdK/-B����?�CD�׋5�1�A����")�g�ŖLy�a���Ida��	�Ƣ5���'5�@)c�<q��'Ҽ�sc@�|�8���G�	r�@aCU�9bl���'Hr�' r�'�剅#���K�G�̟�CD��u���*ä�7e#��z7����$	�4�?�0���<)�������ɹD���࢖� ���JP�?��]i�ņ�w<�u���U�4���I�l�����W4m��`�%�;%q+k�
<�^4B�� ��T�p$�>�4}��n�Op�$�O���P#c�>���n�m"��ⅆ#��ՠ"CH�Z���d�OF��[4�l�3�3��DHĦ]�I���	�*���&�	�2�\5�s�J���"Ȣ���$�A�=�B�4�氀��f�Q�#��<�cݰ������y�I��)�-=_�A��O
�r�CFy���O(���E)��d�Ol�D�M,iq�Φ]y�=@@*��'�����O��`�`�^�<�	џ��	�?ٱ�oHN	�4¢�N��(@�%bR�M�d�&�I���I",G
�Ɏ��-�3=��сdE�6��peFظѼP�elY6`V�a��R���?O���Y�?qŭI�A剕_j�� a�ZX�� E�R�����*�������?	��|����?�)OLL�c��1{�Ho��#�(#��A�Pj@Z�#�O���G��I!#nJ�(��I��M�0�ߪu������o�B�� H�{��פ4�RQNJ�'�I�"�oZ���a�S�? �<0�xIt�E�#���b��'�V�dӔ$���{�)�O��d�O�)�9��ʧ,%BX�Q�N�ю��M]}Zz�B��03� *+O���럐Ii���O��DZԦ睙�:�xe�!9z�(!�/�$neR�شJ���H�K���u�`lqʟ�AT�u�M(f��3�ّ1%O�S�象t'V�f�)͓Hޜ�N�OP���xy���Or���C�I����
R&�K�(�af����Ym>�D�O�D�O�˓]�	�a�!�?����?�D�;Q6���J����!��?�IW\~Rm�>���?A�  ^?1�(����&@-SH��sC W�5ᷧ�ʟT�0�� *�(�pԘA���ź�B����h�!�mN:u�`%��R��TQ4f��w+Z%��'`2�'7,X���x�O��y�iQ�Ff���i��w�lx"â�*B��F1`�Aҁ�'%rpӮ���t~���O�n�-h�I��K�;���7�ZzD�91�#o���ě�$Y\�$fo݅j��̆����A�fr��}��@a�B�k$����n��H���E/bX˓p7b8n����'Vb�'����ݗPL�I$j\ &�H��	$1A1�/���f*0����O��d�O�ɕ�J��S�| �ϛ�|R�U b*��`Ѩ)O��Dh��hF�Od����-L�4�O��ђ
-Cu�X�IЈz�
�H1�֣S���gмk��\�w��Z�'<�mr�\��P��O���K��9S���ui��X(��d�&�&#��?����?�����Dk�P�E��O�|�����ju�(A+
�$A��F�Opdl��H��,?�"Q���49�V�۰B�Y�n�D����B(v�
���m���xr�@��y��9,μA��3����ͬ|2��w�>���SXvd �tR���҂��@�J�y�O@ra���ɄxA��Ń˸vCȥ�"�;zy��D�O��$[�fИ8�?�@ߴ�?��m��<!t/��S��qs���I�	�4.C�8�,94tk'"�Ɵ�S
B����Bt�	��'���s�c@9p�fA��o�	
|��!b��! �����2+O���	" ���B��Gʟ���ݟ��v�ΗL7ʑ���
+��	�4����(�	ty2Z�v)d�a��'���'��tJ �%mX��c��`�&m�"��nM�4�'�b�>i���?�Ġ�F?��
Z.����6^u���V7�"��`��~��w��a<��mZ �ژ��u���y�bL�&g��+ ���tE\�l���x�c�5Q}��R�P��� ��?q��|����?*O�x3ENu�J9�B�L����%�hH���OV�D�����	6.Y8���	�6��be0�O��$.t"� �ğ8)�»�|�	f
	/ߐ-�	�@� `
���A���y����i�@Z������|+pm�0�?aq�'��|��i��'\��'?�TJ�^��'�\S4lC4+�
$�S7\M��mU�1�U���D���?���e>1�	��MϻEt��pf! 2&h3��Q�@ ��Z��?a1�H_?y�F �e�P�'e`|*^w��Ɂ�Q�=$|�`���,����n\!y�0t �'�TAIvR�|#��TqYeb-�?Y�%�(?���f��)d����)��?9��?������
5En��
Ш�Ox�$�O�hR +��[2�	 �	�;\��X;���Ot�R���x�O��D�OԽ;b�O�z� ג��)RB��.��5s���:)0�Ù'���BLγr��VkϿc��Өoq���3`�qRa��
2Y �+V�<����aN��?���?��Iɍ�4�jH~����?Y�y���7ab�]٢.S�+֬���b_� ���?���Oϛ��'{�݉�O�L"���QIӱj%X��(̀An�$P�U�E���$��>�&��Bdݱ(P"��<Y#�08 �}��l�RJ�\����ϚjnU�$]ah�@h��M��Q���'���'��4K�9�b���+e��j O�d1��]�P!�O�<�v=������I�?���;zkW��8�P�)l0
��!���:�M��i��!X74O�X�aQ���i
+ߴ��P�-��X���[}|��e����H�<O�y5�ө�?���J�	��?�$���og�`2D^I�D�r
[�nG޽�	��?���?����?�,O���Ù�Yۺ���J��S��s���#'j��=B��T��ɄX�
�e����Pl�E40�@�2;���a�;TmָcP%�4;���xP��>'H�ɺ{C0�� ��0�����ɜ��!鍔�6�@�R��lc���2y:M��Eş|����(����%?�ݶV�Z�B�@$M �@s#߯�e�I� ����T��hi>��I��M;��Krlϓs�x�@D흴oF>����9%%C�-���yRI�-p��Śu���t�ܿa��Z�)���8~*l`2G�O�W���r0d��Jv0�A�@H�r�Ъ �˓^�rl�{�^�b��'#2�'�))�*�.�Ҕ�η	��a��'v�]��FME�G���������I�?��I�o+4,Y�Í�{Zn�sh�6F�g���Ο�I���ɵ����<���Sǫ2k2&���ɀ�^C❫iO&W���K�%kӐ@!��v��iH�qL�DD�B�:�^�*�Y�->^���Y'�O2X!2q�'���Zc�Ƞ������'�"_���RO�"�	��D��:���E��x+�m���I'�M��!#�p�'�v��?���R��t��=4j�K�؁�?�A]lղ�1DK�]=x1�Q�t�Qd}��!C�U9�"�51�G
�;'��'X����O�`ᒊ��w�j���O(��쟬�듩�|�"��=-?��@M�+*8`	�3�di��B�?���?���py
��'�?�'��y�Z3I�B�Q M�K)|9�-��u*��'���*�'X)�B�W��aD�j��.�?~9X���>yɰ�s���$�@�Of���锸w���O�H^�,��ߖaP�M��'۔|��βR�V!X*�;��! �'�"�'�rQ���A)
�C����ğ0�I>w�F���
&4�T`�ꝰ[���	*�W��	ޟ��Ify��I$3�
��͗L�4$P�Ț�~���j�D
h1�CM��p��P�#���:WP>���M�O��ӣ�T|jLq���CH3�y���y[,S���?��E&�	%�6���?���?��bL���cK�XT�1��K�5�?aDJ�+�(����?�B�i*�AJ���4���ŞMv�8r$��/l��G�	�-Ҹ�Ci�ʦ	�fȑj	�;+�*��'�> ���o}�? �P��J�!}x4@ڒ%�U��"�B�S�剩�?�� �
c������?1���:B-�-�l�S�E�m
�� �I#n�HS*O�1��Zv_���O�����6Y8�1����!,R��S�H�x-�q�̫.��=�'���if\��'�2�!`K�r�dY*��͉2��.t�ص	\h]Թi����3O<m��̡�y�T��	4�?�1�HJ���aC$ ���J��R*���%^��?	��?��?�(O���AE�� �DO�/!����@76�|X�Zb��$�¦=�	^���n �	埀�Ij\H�X��٬w1�A���l�Z,p�
��2����KU>6�I�y���@Ǵ��� ~��ӥ���#�Z�4D�16�\�~���0g�`@��@Ő.�?1��?A�'��q�L~λV]J�"�Ğ l�T#�G�(oN�J��?A��,|�xwJ��|�6g�V�'�M �'G���G�J^p��e���@ğ1�~bF� 8`�*�����#\3G@� ��l�"lFM�,S_�����vnv�1$˒���$��|M(˓4
���?t�8��',��'>��Cǀ7��� ��*gd�A�'S_�X
�4W�]�'��O?p�H5vg�(kU��-�%ZE�9���yy��'i�F���~ �0(�2��'Z��
;n���ҧ��ae��+k�sܴQ:\Ԁ���Ҍ��<�1��c~�
���%¤��k�p������F!:�3Zl���T����4��$ۄ\$��p�F%dر��R̊esc� �<���O�em��TeI0?�%U�T�	D��,�a�Q�BH��MɌk.���4���?)��m���|�%e C�ilxQa=O
�i �Ԁj��<�	�hn( 6�'�N��9'�L��4���#E��`"A��0�HL�K[�;5T�U*4�(�@��ş �I�P�S�_��'v���w7��m�'	kPP�Vf��xm
r�'>�&��~b*M�cM�Y�O�D-� ���Չ�
�TM�1�W�^�� �P f�I4!g�(��5O܌8ı<��'��9
%B^��y��JNr����N [��DP��W��0<)Q�W*p����?��L��W��D>�ak�m�����R�$�'����?I���]��|�hjr#X�h�tM�Э���\�vG��#�<�Ib��4A��U����,�d�$�"�y+op!	�4�0L�ȋ�J@�����OP���O�X�I˰B0Г�,���Or���P�u��Bn�h4ӵɢM/��dV�	���p�O��d�Ѧ���,;C��Ӽk�i�&"�ᘓ��N�<��F��v���%f߃)���	��CT��఻�BxcC@|�hZ�����i��i�vL�"�0����$_��8Q�uj剏�?!t�ÕD&�e���?q���"�I\+.	���_��Z�`v�1d1�BT� p�A�*�6���џ4���?��E/~>�	L�^�
JF�w����L�Y!n���O����O(̪��O�T`0eM ��i�V �`PJ�ِ sT�]�"�K4�	��\ӵ4OܱYҭ�9�?a�
ap��?)"@�f�ȡIFE�4�MR�JL��	��3�?���?q���?/O.�(���/8���۫on8�s	�UW�1�Ld����	�I�l���H��Iڟ�I�W��`F�?c^(K�$��j��D��� �V�j3�I ��ɔ'���h���$x�� ��i�������.#��y�f�1-��8�![�=����vf�ܟ��ş��ӥ>'*	%?�	)X��!@�I`��EkG�d�ژ�I՟��<|2�@�}>Q�	�M��G�f��lU��)�N^7�.����� ��V%�_?��Z%NFD��i>�sC�^ں#�ϙ�y��ވ8T�,�A*I�T���LК0�XIE���X9������
Пd�#�������������1{�% �D��1� I�XxV������'���{WL��u�R�'x2�Ot�,B�-͝'��IH�)��}Pa�Y���d�~}�(y�z�mڦzx��I.Wz͙�3��@ǀ�(Y�%�����iS�K�.�pjA!u���Cw��i��N)����^�����]���C�Jyh9�m�Y��LȜ3����3�'��O�r�'`�I4?��¦A"#^UY�n�n����>�p4��՟ �ٴ�?i�\~�n�>i�i�����I�+h��bjP���R��>m2Ǌ���i$��24��DS'�$L9]�M�Ḷ�y�j5����P ����BPi�'�?�T�'������r���'��O�"%�X>�B�J�";ٺ�scn�U�q�&B�e{������	����SC��S�������W!�-����FƔ�xz�p��аA�i�h7m[Bu�;�|$ɟ��!�@f�)�@�Mm8(������y�g��+G)�Γ~�Œ��{�T8���Hy���O�,�EĘ%�dO�%l��.	����JS <���d�O>�d�O��tY�U���?q��?ad�w��<A��ӫ&O�E�ůJ�?Q�L�x~�>Qļi(46͉�ez���j-�s�K@�6@v�sm���
�U훐�yRD�$=oN�SS�i!��!�T>�cB~�hH!���B���1�B�����P��ۗ:ux���?9��xhi�U�䧾?9��?�C@|8�+�69���(��?6c��%�R@���?q�i�GP���4��� � �|̽�JS�9�\Ӧ��o	�r��O<eх��>�@֝�)4H�N���b�{���ć5úa�� �)j6��Q�߶K~���T�T��&����Q*Ԟ�?i��?��'�Z�3UF�=a�e$E>$�XCI
���dF� �3%�<Y�������|��O�P��(Ј<,�q Ȃy�r���Q�dpٴ!�����G0*_ ��͟�Ҕ�I���\ IZ\�����{S$������DJPE�����S��[�UB P(��&�@8�Mڹ^^$}Sq��&����?	���?!������@�V��O��2��s�D�c��T�>��cA�O�mn�ҟ����;?1Y��ٴ_l��n�*2<p8���7G�d�b2bJ3g�����-��/`2J�1�y�IA>::h���lQ�R"�|b��w[ 	�A(Z;d- ��_g0HV,�b��h���')��'H��)/w��y�Ddh\|���-b�l�q�E#o���'Z�N�7VqƀØOlr�c�����#_��$X�o�&Q"�(A�O����aHC�g��U�Lr�<�c��U�mZ�?)�ЌںS�M-}:BlH2�� j�2`�)�tc��әKt��ɇ� �?Y�3����?I@ML���?Y�)��X:��E�MRpd@���%���0��?i,O��1i�5-����O���韔���A�bq�i���\��1+E��	��$Ӧ	(�4cFVl	�'(��YD#��|2�mH�1�f�'���!�JL�"�A�6�/����F��y�'C�N��	9 5n!.O�!�Nx�"m��	Ӈg�V�`��<��M@	s�1�Iʟ���l�ITyRYw��˓d�,@��Q�J��]P�o��WM"�'A�6��O0�HC�����O����!nxY	�I��^��q J�A���וE�J�&'6��r�4Ox={&oL?�u�4Bo�Ń�'�\��rb�&�T�"*��e�����P""�18�܌!��'�2�'��$��/\��7j�(��C탕nOv�	�b6�Խôa	�n�Q��ܟP���?9��� �U��y�3	9�AZBl�Թ9B� h���'�f���'"(qp�l��ƍ�(��N��e��цe�UZ���۠J�@��au�t�DZ�t�[�9��ʓ��G�?(�bS�'H���W�k_ȡ��L-�L�*�?���?����$�vb[k�M�O���O���P,
���"ĚL�d�Ha	�O�ՒS��|K�O��d�OJ�a��O����O�zh�8�d�+��%c&/M(Ʈ��'NB�ӠAߪ]���)CV���܂}�RG]�(X21Q`��(	�l��>-�L0z0,Zß���ƟlcF�H��d�%?��	�4��)����S�9�u��
*���I�N,� bf��ן�����M��`�z��y�F\�q�ƸY �J�<�$D�ի̖Dl�m;0��+0BH!�v�ئ��L	��i���aH*2^�N�0'@��"�W�g6�����xa�����і	��\ ��ɟ����?���G�+;
d�ڤc�����@@??ꡗ'��X��id��'���O��t��O�b�ǽ�z3���Sϊ%x�؜[US����ӟȣ�A���zP�2����9Ϡ`kѩ�0�v'�A�%�����%p���<�Ҧ�)���ɷs ��'��D�o�|���["ja����5/����� ��?���?���?�,OFT�Ė.-t�d��dHhk�ޱ}n���i�����
���I�S2v���I�l�	�=�<���_�r>��!dۗZ:y#���N����:.*�	70�Ʒ�6D�^�ә��/E�Z!#H�	��!3g�3 (��EB"0=�y������	�?�r��Y@�s���a�4��|H6
B�� ����ߟ���ş@������؟�޴�?�R�M�<��`�!<+n���lړ z���6h�48,H��{������Mϧf䬺^w����78O�Hw٥;��Bô���a��
ΪY��'�����U�Ĉ�F`L�RF@̓lvhP�H�(M���@�L��6�rIDx�E]�v�F=���'��'n��+ă]��|Jt/,jh�+�˟WM����O
�'�6m�Ӧ�CeN��(��+ݓ(��M�:�f�`��[�h)�����,:EL�O�6M8'h��v�h�9O�V(X��	1#�
�%yd��: ��ht�S�Xo��F�T?��K��'��O�b�'��ɝGb>�ۗ��)8�N�t
Ã<���"��U�q-���Iȟ��۴�?��-C~b �>��i����jүUd�ba��ݠ�R�n�^Iڃ錧:!��� /�x��DU�T���1_�M{�a̅�yb.�9Hъ����%�`��p@���ɛ�?�q�,����?��r��7��I�o~$��I>7�1�M,O�X!�3~���D�O��D����6��D�٦�!8@���X$Ov4pp�eш>����۴M&�S)�~��Q�R�&��O�f�Y����%��$)i���:�&L�PP�a*u�C2���	�b�<YE5O����Ţ<	C�'�.M��È�y�,��>�7��(u�]��AP>�0<�5�� k�C��p������@��;�:�A�0�T����M�41��%?q�_�4��џ<�/��<���
YPy�!�f�m{W���g��y�4O6�o�
�:��7MV:f F�'K��͓���9�D�.d�ɨ3��6G����h�'��;��˓����'���'@(a�'�N3zU@���0�����'vrX�׀�]c�'->7m�Ol�7���]"F4��Z�)�P�ıc��&� %��Ijr��I;��qq��������yr'�,6B���;F>T�Q�y����h�I�(��鎺�(�6���Q�G�|M3S�'��'��ěs��`� h�����3X�!���}y��>���`�'�b�'����˱���'��,��S�^��Ro��L���̨>	���?�&HUS?�2�W8Qq��cs���tE��3G���bQ7r��:�4W�|5:�'X�<����<2�Ӟ��[�����7����ɕj�� �"[:Oh�|DJ5LO�5����Y5���Y&01ʔ��T�6D�\i���B��$�ۦ��	�[N��6e�	'�Mc$�i�0A���(��d���E[qm�0��4�h]��)"�'�@@p@�̺oZ0n��O������8��J\8�0S�P5*��x��g�&s ��O����~��]Z��y�̃ /%RL/IKZ5�h�����[���?!�r͆����K�|r��y@���'��i�'ɀɻ#_'V�НAC
;�\���,��~r�Q�����i��$�4kN�NZ�u�4Y�	�5 �d!B"�i
r��OY�T/����" �$�C3>ʓ5@�A�I�\)�yR+Ai�%�rmU!7A
�i�G��O�X�WF�5}�����O��D���C�I+?_��bbjO�m���f�#:�����d���hݴ1����3Ď$�pe~>�{s�C9'�h�h�l�qZ��#)9 <�+��%BB��<�S�r���I� ����'��k��C\��k	>?H:��O���Ad�<,<���O�i�O\��<ab+�2	٘�B�D�*&����/�T>��	!�S7�?��p�F�'�ڕ��O�'�V��H�d�(i۱E� 0F�"k�.7͗@�J��RĆ^_���:Ovݳdl��u�@�
�̓��I��H�S�l��tÍ�n5*��I�?9�(�L��Z��?��z$�,��I���n�h�U����^݊ek��"����O����OL�)�P��O��nz�-�0k(o�	����)RP탁E�*�M½i�l1�=O ���O�-���.2����XL� f�"�m��}��Y��_qlNp��6O�tj�cT��?٧��o�I0�?Q6B���Q"��b*a�4��53N49�a�7g�p"��?Q��?Q)Of��Q �#$d���O(�	 VD��@�H�/Z8t|�s�L�}/����0{�I����ݴ�l9A�'���,Q�I��A��d���Ý"-��̓V=t�P$��t8�!���}�4.���?q㛑E�&1hc��	b�j�X�OU�h��O$���O��!�4L���l�D�O(��ɭ&��������.�����>/\x�K�O��黎�	���Ӽ{�BW
6P�	P� 9wi�-ôJ��I�8q2KU��?a���?��a�Zw��[�1O��/��uߴ?�������,���hr��s�����(����DVɟ@��H�#swx���������?QsG�Y津�HP�c�b]@�c����',Yi@��3"�'e��O���	̟:!ɰ���*�~ x�Ǌ^��ö�P}��'��`��~�āYh�OT���@�E�R��C���I�2$�Y�k㛆�[!_�݅by�8�'(]�%_�Z���
�@@�A;�b�k��B�V�ӧ�(�� ����?���?A����U�R��l����O�:7�17���kjG�����B��O�=o���x�Ƭ<?�E\�x��4u�F�Ѕl�f�@��K F� �ujK&n� �rBl�V�м �$C�"�N'�d���W��������wݖ��R"
�X��"��b�N��F/� B$"(���'oB�'���`1Y���yw�(=��`��-e�zp�r�ў���'$B,N�_��܂�O8Rdlӊ�D-��H�I7��I�ĵ
´\�f�Tj� �S�O�����	�NH�O�l婖��𼲁 e��r�=�T1+��ө%6�9��B��Ij~��w8O���T��<��'��٫�n�<'�'��n�P%J�J �OS��5�'�_���'��ɌY��<�6���I�� ��V�l����a���B�S@�U҄�=?A�P����ӟ@FE����o�6P��2z�A3֍�w28(�æɋ9�N 
��0�6�L4I���
��0Oa"���<�SFܹ%>�<ku��>;���F��]Obn�9B�
�av�'��O�r�'�	W�t!��~�:"D�c�^��$V�fA���c޴�?�S�GQ~��>�������k
�%��ȴ���{'�����(������ q��`d��<��H�*)��}�(%k��d�Ժ���;�&ճ ��J-�q��n�O��	�_+B��3NUٟh�Iğh���#B̕O�>AJ�b�3%lܻՉp,��nڥ)����'���'��t�[���C¦�/����]	#
�'�Φ��y�	���8A���K7(E�_���=UMp���*��k⨘�8�Fع��G��¡��y�ϓ4A���0U@L )O.�I�V�HP��	C����D�7~�6�#w��Gz�$���ɟ`�	����	Vy�
։5���6�'_��'���8w�%a?�S�˄�L� ���'�P3�O<-�'���'�Lܻ�'YN!��.@�M���e�R0[��	sR �$Xٰ͓^��{�ː��ٛ�)]b��㗮�?	�B.p{��X1C[�;�d1'+�},�Ej �O����O:��tY������O��d����ׯ�6CF��ǘ�4
��*	�`$�D,�O�������o�j�Ӽc�-x%�����	:����#�"&&��n��v�'t�%a'���)�Cf��Q�ƙM�i>�8֯�R��]��.X�:�%�`�G���I��?1á҈�������?���$h�<� ��Ra8�1� ��<c�jq.O�ѱg��Rӄ���O��$��&��3���d��V���I�yj�ͱ1R8�d�'6�6m�ܦM� ����s��/�	SW
�B��S�#F6H�F!
	in�[U���uF��<	��"�	�E��'�����-�=BGc��V?�XY%�A96����Ý��h�D�OJ��O��Ĥ<����I�^��Oz��FK0<U,}c��=K�A��Lj���'4�)�Oꅕ'���i4&�h�� �n��ʍ��~ p�*�� ��X�b��	�p��'�&p2Čֺoa���O����C!�b0�*&�*-+��ρm�P4{'F�����OT����� "��)�9��Ec$X8nY<)�U�9$,��3�i�O����O��D!	�nK���O�o՟��+~���ǧ��(�p)�f�2X��a�(��|C�=ϓk��&���M�'rzdZXw�����:O�S�牴f	��aFԚ

<���
�D[���FA�CX��c��#�֝�@�@�D�O���!^V�h���Fx0%������O�";P��B��?y���?��'Ta�h�AI
�,"ʠꦢ�}��K���]~+�>I��?�2�o?1�C�:.��*QᲽ8��(~�	s��,v�¨�P*�.�(�lZ�e�����?� �%x�Ԇ�`y���A�&tK�S�~z�"��M��l�|a3	�O��4�8��O8˓H"|�+��P�e{KG&-�樃!N�
ɐ�����l�ɢ�M+��H����'�`꓈?�tLA��jṓ�ț[)�I��ٿ�?	@(�uȺ|�f^�W��͓��q�fh�7�� ��I3jc<�#.�ݘm"���:%�>�$^�Л��V.h��I��l�	�?1;"@�w��ӔL)��Ѷ��^x�l1�`�=��
�AE�L���'2�O�*(�Osby��.����d�	�,�J�f�K2���O2x�7�O6	i�l]�G�R�O�(�����r1�c̈́%�L��f�cZ<I"�lUHb��I,Pb��"�5O� �'�<�1�'�q� GO ����'�&M�F��� 	29��'��'9��&@�lB����	̟�:� փR_�]���5*g�}RpA�8ّf�p�I���čΦݩߴoUl�Q��ti����I�lhbӄ� �8��������I�Y�h�4�_঑D!O�<A^wK<E:�'����"�,<BL�1el�t�>9��Ҳ$�"�d�O
�dH�GR���GE>���O.�4���Zw�R����`��=A@^�@���O��PE���^d����Op�nZ��0�x���i��h�F��u#L5X��5hc �J��F�DL��%�-�M#�D�7�x��\wh��rѯ�O�����*�u�4XlĊ��	����@5D�ІK����KJ�l����H���?M��HN�q�� !�6B�|��&<h�6�'�E�1�/�b�'���OrNi۟O�B!T%`���a���G�4���� 7yT��?a�4����Vh(���(�#`�? > �e�j�z�(��]�`y��s�ج�p�r�,ˆfH�/��_b�^�r呚C�T��fܡJƔ��E�4NU~l(�k�#\2�'=�'��W�0�â�4t�����	J^Hx�	�	$�49����8sgd����M��}6z�'^�m7�6�|�NT�6�[2��iBP�]p�Z����֌�HI�^�ȕ:�3O��F��u�4����*��i�ݧ(�Y`"I��$y�JԀ�3%D�&
 �I۟d���?5��X^�s�qR��کCA�i$�1n�A�O
某�I۟ȃT�_�)�F�S�$0�4�?A���<��_:(裡dW��k�J��0�"A���5rGިDm\7=�R	9r�wݹ�E��<9��E��IsB�f(�3M�#DH�Q�z�$+��Qy,�O84y��y���O �$����M����c,BP(��H�j��D�O6ʓ:�. C�%��?����?q�'H��M��I�"E��tX�PZB�*���x~bj�>)���?A��i?��ܱ5l|�( XD)z�bX5TZ�,�L�ꈲ�AT�fZ�}m�42�ry��?u���k�@h1�Ey"�L-/|#Vc�pe�|���_R���;��ɛ�F�O��4��d�O�ʓ+�̙hI>)k�}�%���p�|H�񢐎A�ݱ���?�i?��I����]y}��'7V<�%A78\!Bkf�ȳG��A��&�A��Yl�n8�r9����'��iô�:A2O&��@o��Q�����H�*���'�$�IM��Y��O�$�O:��Ϩba>�'kf*�ر�P�*$5�V��R@L8����keVm���?A���$l�S��li��nS9+j��J��Єo"��#�	h���D�O
I(��O�h�
c��O�8��S��̀X��'~����UH"l�M�`9��:e�HI�4OD�#q�<y�'5��� _K�G�r4�R&<45`�@#D�l�2�'w"�'#剤:�8-�¢������럴��bY���勅5�R���aWٟ�CP�$?�`U�D�	ɟ0X#���jp �Lw�iB�@�a+�m8��U�'���3=O� 2��މ.�D6��k"�'j�H`͓NN�y��ϓ�B$|��@<_� ��̄ ���'��Z;k�~�����'���'���s햑r���_)�8���'����vk�G���'p�6��O��ƛ��]6e�Q��a߱X�b��	[z{�d��U�Ν�ݴv\���ET��u7��S-��=d����[w:��"-� KT����(�Z���!d��'���D� $���tm�OH�$�O��鎴rU���"ϝ:%!�!�2�8��t��<��^6��\����?���r��H�|R�t�L)A(�=ZN!H�J��k�+�]���IҟT��#���cv� ~���1\6Z�i�$=���G��M���x�\¦͹��T�<��o�!���I/q͖'xF�D�oZ�H{ѬظT�ې��B) 2�P����O^�d�O���<���X"q�j]��]-������b�\��I	����qC���'�Љ��O!�'��7M���j�
Lc%���l�
_!
@yD!eC&��A�4�l,�uFE�<9���?�F�]����$Y>���;&��-� �m_�p0�ɼ����I���"���?����2@f����缛�Α/}걡�,ϩ혥ju.ݖ�?���?9j� ���O��7��O�-��0O��I3o��R��I^�4L����G�d�n�3CSԦ�ӵUn��;��@r�'Gl���L9yj��D.ɛ=`�=��� ƌ�	-
�6�Q/O�e�I��B��4
˟�I՟d�աŉ!G,Ms�C��1�\ii���Iry�&��W�r�B��'���'[�T.��AMz���<[�:��Mօ��Ol�'�³ixX;�'���r"���|ʳD�^h�s�"��8�(����V>> 7��\���ҧ���O�Z0�'0���!S����nC�%� �b�-�_9�`�¨D!�?1W�C�S+��@��?�'�?a���ŨW��q�&�[�*I�M�!��C<J�@�l�����O�4mȟ��v�$?�`T�\�޴"ph�{D�A)�x`��V�lQ�)�i������ޛ=_�y[�%�y�苉>7*����9��^�<���)(�N}v�R'z�aH�HT��d��!A��8�]��?���?���6�2Q�/���hB�uxT�c����w�� �Dd�e�UiT��O���O�����@���Obnzޥ��J
o�������+�-�bY�MK��ir:8��'�}�FK�s�Ԯ�R��.N,:S~����7B�s��¯|lM��k�l�`��GO�D�-�^ʓ���>�#�'g�A���׿n�2]�0�\�f��e�'r�'rX���w� @)J�	��4���(���W����'�>F	f���9Q�t�K���ٟ������I�"��5����Cm��r/�4p��I#",��D٨� �bDIbӠ5��.�|B��U�<�D�B#7,T7��W�ĥQ��֟O��yh�'�'�h(Sd�R!y�O���y�B�mvB]2!J��M�da�S&"�ݭQ ѐ�'�r$vӎ�FR��iޝ#tk�
me�ek�d-U-X��!�߹4m��ksaA֟�Z�`�#V�ŭ�d��]��'�f<S��ɺo�6j:�A��cݹ\�a�u� .���-�~yr��O�YҊ.�����O.�D�h��s*��zF��f/�.T:�@!�c���XBd!K每��?����?Y��ט%�O}�@7�ܽ2ԑ�'\�2v� ��	��`��c���	u�v�CF�?� �P9%���ԨL�fJbؓo_'���mZ3�Hh�zPh�Є}���2J�ky��O���R��>qF��0+�""*5�Gh��VU�i
���O\�D�O����O�˓Y��`�r�P�?���İ ��ܛ4L�GT��b��?��i���\����Id}��'qb�ͥ
��]�E%K�*`t�E�I5�t� �j�j��+��ד�yB�� ��I��F��TH`f�|���w�}АnX:c�~qh`�"�����>8�,�q��'72�'��ċ�����y��
X�0����,��1�D�O;���'d2Ѐ%:�j�����`޴�?qe��<�0\�Hj]�B'M�)����O� ���ds�OB����|-9P��|�Jؠaj�%2���tr�*E���!�h�%a�<ઽ��(P�kʵj1�\<U��/پE�*�ۗ"Y����̒�Y����H��.��ɓT��a��96HP���H1͕#wѰ :t
ԣA�xA@�Ʉ�0��&NMn�d[�&Z�A;5&�Ԏ=���W#ku�=s⥞5Pkp8#�MY�z�^}*��6-B�)����6�̵ɦjӪxm�3c� :�����/<2�����e����'J�r-s���f� i��G֧k�1$��5)T�(ʆ���II�q%^�@()ł�'<p�``1h��\o����	�|\ڰ�@ �-�4�6��K��8�i��'���O긨��O���"pm7�����Y�~B� ����|Fy"�иG`�<� �21A0���ӭ�M/O��hF�צ��������^}�'���p�@�^�4J��a��m1%�ǌ������=�&E�ZۈB��:D�D��e
���M���?q����T��:���O�#G��@'�=��M�s`PɪԪ�����"�'�r�$\�x����{�*�Q�Y0e�6��Oz�D�O P����@yBhO��?��l
�l!�-	�� tL0l�C��HZ2����O����O@PC7e@�<?��CB@>�f�i��ަ��	�� �/O:I!�'��.�����v�c5/Q�Y�B�i��(LY�hr��I�����d�'�N�
A�*8x\�`���x:��C�U�V|xʓ���I��p9cD,��Ox<34ɂ0�U���� ;SJ>�I�H�	� �'�p��$~>�&��(��@гY`�S5!�O�s��'��K'����D���	�<q�N)�Ac�
�z��Y���듕?���?i-O�h��A�ӲS�H�If�hzԊ��Ƕ\�T���4�?�q�z?�2DOk~ʟ�_�R�x`��=h�-3�B���l�ǟ(��qy����(�f�(�������.�#!
e�/ҳ8��| ��Z+]X�$G����C���d�/t�8$�p/L(,�.|ht@E���^�d��*�M@_?y�I�?a:(O��Q���#���7n�*��	�lk��	'rva{b�O!\aL�� �Z�T�H�b�:�M��W�3��'���''��J�<��U����5�Щ �ٗ\�Pw�=Z��ً�?	�a-�O�R�\U�����O1)�,�a��u�~enZ���	���㡁���$,>�'W��Z޴S�JE����q^&P���	#	�A���ȟ��IꟐ� �ԓ;�����Ō)� ��Ǝ�Ms�Z��h��_��x��{���	6%���kL
m~�Y0a�!N|T'�K���P�
c�8�I��0��xy�ǜ�I���qd#J"*o��cG'�5���h��>Q��]�<q��=����?���ßDQ���/���Y��@�j�~����<j�,�&�4������\y�ŷm��Sd�T�A�Z�g�у�ɀ��6͚sE���Op��G�O�T�'�B�N���J+zC("��B'Gh���'/R���?���?�*O2�����M�t�'BR�]�r�he��D��Z��4�l�h��"O��=�R�'�p�)��$K��De��k,���N�H��'O�U��`p,ߵ����O����>(�'(+�	��n:=�TC1H	m_��X R�':��!��'x�'IB�]�,NX2���'!�=�W,Lj7��<A��9��V�')��'��$��>a���-x3R�[���5E����0�D�	������?Qơ�8��'��1�M|J"�0��試�R/2���-���)B�  ��M���?����B�W�����b���SC��l�ꭨ�eG�Z��	p�eG��M#�E�O�'��YQ�y��'���cw
�D/��j$V�[ ` �i���d�O��DU�S�"��&-���?�jZ���C �L�U�Uh�04=p!�4J4�	Z�Ι&����͟�I ,Q6����b�`�����W��ܣܴ�?���ͪ����8���՟x(g够����I�ȁ"cX�Cgo��b�h5��Y�T��T{�I����I���'^t�5��#j#���1��(��M����kk|�[F�9͓�?A�/�Z?���� ��%f�0'��׎p��<�yP�Kϟ�'dB�'%�[���`)�����C�^�Z���+"	���c���Ms#���<q��F���?	��˟���L�w?�A,3,�lK')�V39�GF�H}r�'3R�'S剫5�܅�I|��߅l`�j��i-��s��� ���'H�'Ƅ� *O��Ol�T?�B�'A,�� A�q���&t���D�O �H�[C�����'�\c��u{�^v遴bR�d�|�{T	��aGo�<Q�����d�O�s��]�~We��C�9F��2@�.��7ͪ<�rI]�`��j�~r��J�Q�rE�� f�Sʕ�Z@�wꙵ;Z�˓Vrtz��?��yʟ�������u����tܻ�F��Mk�cIӛ�'���'����<�P�x>�K��>pu��r�ML�t2=�FH�M��J)�?A���S��'6��e} ID\=r�^��&IW�27-�O���O� �S�fy�c��|�vѐ�o�uQ�4�׃֊J�N��t)�*.
7��Ox�O ��<���?a�����,��h$#Cܤ��`�O����"o�=�'Q��ϧ�?��#Z�D֎��p��>J
-[���8e�O���$��|��?���*�Ь����8_TP��"j�?l��9K(OH��O2�ɷ(��OY�ٟ$x��Cu�buA�٣)��وb�iA�u��y�'q�I�a�T�⢕�r��HQ+E�H:Iӧ(�Ϧ�j#Fܟ�͓Y������$�|2�T��M��N�;��Y˲.h.i�@�>����?�����ESr�m%>����x@u#Wi�3�<����M��o�%�-zH����4�'��Ԅ�'CJ�2h���!H/pw�T���i��U���ɞ|�$��O�r�'��\c���Isڣ]�e��� ����*���Y��O���d	�K��u���6$�QP�lɨ~�dĈ�M�.O��ӓ$�צe���,�$��"q�'�� *='�.��͚`싩 x��'Ք��¾H�����O�s���=�Bf�7�d�ӅM�!6�$��j�@�1��O0���O������O��Χ2;4���7a�Թ�E�J3Z��D�'hF}�ɗb���h�I��mj|��D�P��,æu�	ɟ�	�yt��'>&�O���G��M㲭��i:�&��N'
�C0%E�Q$�XH|���?��jD�A�FD	+?���Vĺ0ži���ծI4�=T"�S�,�Xk�d�%9|�X7I�B���g�4M�7ͣ<a�����O��D�O���T�#�C�K��#�DP�Rzx�"'� v=�ID�N���O޽S&�?���u��؀b�̐�q�Ηf��颢Ƈ�Mk�����Ol���O˓Z� �?���kwf�&�x/iO
T���'��]���?�V�`?��Gy�O�̒2Ԡ��!� i�Nx{�ÜK��ON��<���90�A�,�F��4"�j�a6囲DG�e�Ɔ�,�n�<�"������O�˧�xD&��@���,_��@�h�c���v�<�$�<���Z����.�,���O<���&mc��N~i���D�[`��y"Ll?ɇ������u����O��L�A�T���H�Q�p�PD�xě&X�p�����Mk��?����ET�JJ�JI�A�f�eb�pq��
#����ݟ���Kf���INy2��2��'W�6ػP��D�^��&���`n�&?����4�?���?	��">�I�4#��	{eP=��"��l� ��܉۴M/��'��	�u&�c>9�	�u��@����S�dAY�V_ ��4�?����?�a.�
!V�	��4��ןDQ�Ca��Ly�ϸ��g ϖ n��$�i�RS��X��j��'�?���?q�M���#eO�"麉���<H����'�j�eL�>�����<���jn̓���+���
wȕ�~�f��ĉ|�m�'���{�O���x>�D�O�ʓ~�`��0�#'���eA�%"��8-Is��I�w�D�ٟ�#�Cr���Sџ��I�(䖕��^�;h��3�+4Ѿl(a�{�h�	ȟ\��ȟ���Fy�@h�L��ߴY���̸U���d�<(��7�ڜ}���O���s4O����Oj��_/r�ě�hl���EU�G��l!4��9�l͟D�Iߟ �Iay�,S�(����?���[��q�͔y^H���,��f�'�āٝ'<!�s�'��Ҥ�y��'5B��'59x���!Y�8��x�Eo�)T7�O����<�Rf̝h������	�?��M̴y���UkX#��:ҥӚ;V�U�������il���'.�&r޽���϶�h���Bn2ʠ�UadӴ˓O`N �g�iB�'r�O
��m��lP�;`�ɖ�ŷ'_p�X��
��?���yǰ��'*剶s'��>�S�OذWL*����-K^�ٓ�i�V�9��i�V��O���.1�'[J���'Q�g-S�5����$�aZB�Ѣt��ڪ���<���}̧�?���ڱs��W���ҕ��G��m����	�PC������Ğ�H���Or�Xf�i� tQ��T�������^�1E�}�}����'���'�E0T�b K"{�h:���g�6��O0�)�iPU}¦��y��'�����'m�\c�؝�F�F��|���6[�rD9�O>E����@��ǟ��I�h�'DjMp���BC.��lE7\�h�v��+\���c����?��G�<1���?9��)5x�q�۟e24��� �$KY��ض��<Q��?y���?�+��ܭ`f`�'�l�dj��$��a#� ��o�/g�P��ܟ�Xb�a������������	�=l���̷`�`z���#�f5�O����OX���<� M�;8l����Ā�?*��IӆJ-x�]E�Z>�M��� ���k7v�����?�c���<���?�@%�������"1?D���bRQ���'�2V�ܐsB�6��i�Ol�d��F<B��Yw}p֋�B6��9&-��/��d��ź���Op��4O���<Q�?�|a���D�x�	���gY���g�i��
]�D��4�?)��?���tY�I;L9�%(��A4Os"P��� �B���@��3[Ɉ�����1�Og��z2�F����M��1X}��4'F.ix��i���'^��Ow�+� �ΓNO���gE�����[�:����i����	�1ON���>,<:�JX"#	���� ݳ{��in�ʟ(�I��P��)���D�!N��ON���i/���@G�"]�|2�*�+"����ݴ��F/��S���'�"�'-2����J�<$I�Q�ʾS��<*��������_��Y�'=.�����?�f�DM�\c$���C�YuD�S2E�*�~�:�O��i��d�O����OJʓC!2@���X�<��"��,
S��K�d�u�I�u��O��Z�?U�I�4zsM�N~R Z��'pH}9�I�����Icy��'K��'��	�E���O�X�I�+@�\�ᅔ�_�l��1������h0�#���)�O���D�N2�};��(.d�p�$ d����'�B�'r\���V���ħG߮<�Ÿ{d�$0�8tm�`���icbΞ��~bM��?��=��X�>��իm\>���e�@��l7��O����<Q�*H "��O���O�^�W��!�����E�{bd��F/1�~"�H4�?��)��ѣ����z��G'Dt�+�\�B#��[�"~���X��9T�߃�MC�_?�	�?݃,O���cO�*���� ;K��t
ܺW���'��ѓ��'��'
H�M|J�e���P�tÑ)?����F�U�6�K��M���?����B]���72O^��A�
���C���g~qAF���U�ba�&��9	.�����8 B�4�HU�IS9�.yk����M{��?��r�B�w_�L�0�O
�D�4&ƛ� @\I4���8g@<��l�)0�T�;A�D�-�1O����Oz�єg�xU����D�\�U�ݭ#Yo�H����*��ޢ(�2�'�ȩ�ϟk쐇=m\Q�FJ�vM`�)�*�6N��I�&�L��IXy��'�B�'`�!R��i[u �*� a��o۹M�@�6a����ͬ��'3��ɟ���O.���O�~�3����¤�1WD�d�<1���?�����Ô ���'|Ū�04�ZG� ��S+&��I�p͢�$�OXF�O��'`B�Y��y"ME-|�fH��
��$5��uN��?q���?y*O��J�`Gd⓵J����9{��a)$��,�x S۴�?�G��<�e̐��?1�+U�Қ��I�}�����d�k�h���̀+!�6�O �D�<�d�� c�O�b�O��t/o��Y2�@�diĤ����n��U��-	� �����{�4%�pk�w���%�î3�0�;�K��v=�۴��d�:�N�l����I�O ��KJy�&�,ROt� �nY �ҧ�/*~�q(���?)bQ��?�J>�!��SⓍ90���JTBh�6c�J<7-��B��o�ݟ��Iǟ��+��I7��t���S��l��R:0@>`K�h��	����˫g[���i�O}9��H�G�<���?1����3
�ϦU��矸�I"�4a�)O����OT��K��M�TϘ�W$ɱ��XmA�d�̦i�?� ��d�'-��O��q��F*9����)w��h��iG�(R�ɬx:��S��e⧟��	�5�TE:1��'/8�g+Dsh� $�Ћc )?���?9���H�;t� ��Ь\Zt)���(O��$JyRH���?�A~��O�"�'2b��Aj
h~�1B�L���- 0�����'�b�'��V���3�ֆ��TL4Ö��wHݩ'5��ѳF��?i��ޟ�I�;d�������O4��P�<��Y$O����G�[��y�ͥ<	���� �㞢|
�U�~�Dy��s�hP�OSL�<�$��hE4���䏺]<n���D�_?���Ϥ$z��� ��|�q/ΰ(��b(��1a����B��$5�p��F�s�y��D�!:(�<�3�K�5Uc�z��ܰ� ��$VK�5��t������L�2�j P�����8s�z�"��nP�Ug\F�*�T�_�LI2�9�nI:e�n��fC�$IeB�'�����n�z�h��D�)�,��A3+9�H��ԫ2�F9�p�x}��sɂAU̅U��'�X�S� K0�2�҂+H6�x��K\҈���ua�է��B-��9+�c�a�:e���G j�B7�'b������OZ}3nP;A.�<7*˾n ��80"Ox��TE͌9���r�� Y�tXR��x�q�K�8��?��-ӺZ�F�j沽�π-?_����?q� �1q���?Y��?yr��?�R-��=dH��㍏bq�1[S���â��G|�� ��yLvQi�'��-3F�R�
�R�ͦw�hH*�'~�D�����
v�J�e>O��U��y��,�|�d�7�O�(8A�'b�	@y¯�i�\�6EO�/j�<���O��?��;O:���ۘ���E��A(N�a'N�d����z�T�'����Ыnv� �q� /f���!�<b���B`�'h�'BR�Y�w�]���'!��'Xӊs���:�t��a�FZ�\�mF�Wz�`�Jt؞�ѷm9#��Ɉ�@�������ˌ�-���*��FУ
ۓ{"���Iğ�	UkS�	[�ԣr,2U�@y`� �R�'Lџ��5�R�}"����9)
u�W�7�?�Y����?-���kN�f�}��Iw�tTOh�P�'ܨ!����y�'!�@b��3"�2[��3�&g@M�ę�4����I�� �D�ڀA��0!'M:��԰+$��)G3�a��L(
CL��gnޢj�Q�l�5�2p(��7h����O��ДC�{ȍ��-ѫi%�$����2b���'I�8y!#@2ue
 ��Y84(u<O���ܣsͰu�H|�܉R�DD9��I��HO�S�.gJ�
�$jO�!x#J�ʓ*��8��M�B��7
Q�<�����MV����O���D3T0b�W�V	���q6Ø1	nt:F� .����a���O���HV�����Oh��a�%vR)�$j#��[��8fn��3b�;X����O?��)y�� )P���7�±�C�' c������O,�d:?%?�'�Hi�V/j�>`Jp��[.zA��&&D�x8P@Ԫ�P�U �?P�T�H�$#�DF�<Qf��\��'���r�����P����ŒOe�����'��BZ"1�p��@�'���'?��ֵ{oh�r�'�(8:A$�3������]׾���'.ByQ�?ɨ%��J�9d ���f�[{�l��w%�����aJjDQ���b��A��w$�I#$�v�$!|O~��E�6hW<���N�4&.�����'�(�	�y#,4 ��P�S��X�+ףz�\`�;��?�G{b���|����熏rHH���8>i!�Ě��f����wg.cH		Y!��(\Z�Y3/M)��Ȋ �sU!�$�?��L�©�|�V�"��[:<C!�� ����K�VMz0�qJ�l�jr"OL؈�I"R�v�QdW�$�-�"O h�R ӌ	=6��E�2O
8�5"O�)���<I�	�@'Z�T��"O��KPh9��q�+��)jq��"O䀩e�Zo�pu����Xvȩ"O!K2�/ki��r��50�1��"Ot5(�c�[�@q�¤�[���&"O:ܛ�'�#;V��F*QF�Ҡ"Ot���ܕK�
H	�՞K���!"O���%5	���B����3@"O��S��*��a#��v����S"O<���S�}�$x��nݗ	r���"OU�dԩfB,#�-�+`���T"Od$H6"�S�؈�1lA�D�}a"Ox����!��,)�kNM1�DR�"OBa���5yQt��L�i'2PI&"O�*r�<]yV���j90�"Of���Ժ:C��E��9%�i:�"O��iA}�NQu�äB�U!�"O�����I���!�#3�,h�"O2-�1�̎Ub��A��J�"O�@��BĒK�u��k[�sm��["O�HE��@jTx *� ;NJZS"O��;Њ�V��Y� $�0B,��CQ"O"�1N�Qt�45a=#%�t"O<�ԈY(�-�� �PJ�z�"O���M�tv�p��MTpf��HT"O4�0j��r���/սy0�]�"Oj�B�i�g��p9m M��6"O\��/�(�����k2"� 3"O.��f4jPu�E�O�b���q�ɇ�������*��c>!2��P]n�{@�0rXFlqrm,D�  K�ʀ�j@�	�@"0��)k��z Y����H�"?E�ԅ@�5{��C���.�5JՉ�#�yr��,%f����=U�2hB�nN���$5��E��ܞ>gaxR䊹U�J,P3��K���a���0?q���&_܍R��X/Nڢ1��Ҝ"�[R�I%1��Ն�(ۄ��6�S�\5s�̏�Z+� F|�e�20��]*�J��OC���U��$z� �l�-J�2�b�'����w�0Jl��	�FX��0�'�^ �D�L�d`PP �O?9A�ߑ^���kɵ[񈳃)D���vg��'��X�1\5.��S��&?��c�nT��q'��O����ꎢAN���S��Z?�p��2�O�(2�	�PƵ����9hY�fh�-�(�rj])\!�$|�J�1�cU�$���ã�'en�#�P+7�h���:�S�9�t��#�*$:Z��r��w�B�I�DJ\�@#G�V��@���^�2��ɧ<b�)���[���S�Ov�5"F�G�^eҲM�t�|90�'$,e�a�E�W0����Z�y喍#�OpĹ�I�|��[��'�F��#F H@�#��zQdy`�,�,���Bݪv�%0�dUR�Ĉz��#w��(�]@<9e �'}��*h΢J���GQJ�<I����B�I�kB�A]�X�u�D�<�'E�-��t`e�109��E�H�<��i̾n [�JU)(NZ	��ISD�<%�f%ΤYWE]�wj�A�Dz�<��'�[���+�!m[2Ha"n�w�<a�
A�GDR`��� K,:yyrLn�<�цحu��`��c�x���dd�h�<�W�J�T�N`0�D���|P`�i�<��I�afx�5�Fb���]�<	�Ϙ�\ɉ ��t������[�<��K�$.������!Vl�a�dY�<� H|:�GľQ�X�#�]�Zo�HU"OV�JG�OJ��3`a|�#"O�ѺWd�EJ�gd\^z���0"O�I����4���{�42�"O�g�H0 F���JّR��a3"O��*_7nћS��S2T�A���y�,U�D���Z���Q�D1)��y��G{�X )�D�(�
7dV��y���0�D��q�П9,F�٦ ��y�ܖ\ĈȗO�*S����A��yB.Q�1�*��
�H��;��R>�y�q��4(B.� B�h�����y�-�	e�����E
fڢj�C�?�y"hMT/� �aZ[&q0�@��yR[�<��@��_U�� "�����y򀜚\����F}��2��2�y�C_�
�`{���r1.P�(^�y���'�=����sHa9��(�y�.�'N�����p��4���&�y"���}�b|Y� � F@z ��ybH�(qil�!��T>0r�ۗ���y�I��x F �%�@���F��y*�3a���h����t�V����d�J��>E�Ԉ�>Tp(�+_��p���fI��y� ��4)N%Jq�% ���x�`ځ����8R`;,O��{�G�D��QF��4F"���'e��;1���$�b��
c�H�R(b�h���vt���cZi�����K!+ǼF"◌ma,��~���!k��P���Yd�d�Yx�<�W��8@��JƫЄY{���*�ry+�Fv��=E�d,R��! #b�Ŧ|8��8�y�*��4�H�(�\� )*�Ц+��MS+�y�$D��de��I%����҄�-1!���f*]�o?��$��_\�	�>B��G,	$5,�b�)�(����B"t�!�d��<3~�1�ĿIr�Β7[qO*��
�mӌ��uCߪ},�c?���LU�g�"U��dč8z�+�F(D�X�#� b8�M1!OC+������z�"���4Sr4���4: f5G��OD HC��]$���q!N�Euh�S�"O���C܌v���	�m�n8�+��yl��*d/:����&<OF`R�J���5��O�L׆,��'^���i�+ÖpI1
��
�x������ip�Ζ^n� `�O��+᫚�%kLL��/��s���E%�q���R>�8Y���d�'m<8��48�ZM&c�'p� ݇��O�<9��eƓ*�4���ӥ����(�f=��A
Q�8\�5�L ʾ�G��O�̐W���X�X�0�e{������,9�����j�+��<�'����LRAGG;�⌸Vޓ:rй�5!�U�t��u >O�T���[,W|r���暍 M�! w0O��p�/Ǌ_��
֜��3?Y���!iUlu��D�0���6�<���VM��C�IIC�c�U����A���"a�'�TȘK�H��+/��4g�/"�F70���8�MW$m\`=�7J�<r����'��ʆ'�)/k6-K�F�!B�(�9A$�GYZ%2�O�@)�)b�\9��"��u�$C'���O����ٗi@ �BK�.��P���I?SC�0�6�`�(aK�=O2�I�#cz���˒?j
e"�)�#�86�W�8?,��@b�<p˓ZZ�q�̲M�d�kmZ$z�6�ϓ_��-ـAV�Q�D�sf�OZGzZw�n1���c�4�� 2�DAP�'�Pb��0R
R��N�;�:j�E��!�2<���g��|��t
�2������T+P|U2Ac��o�n�Q�'��)�<A~�ڵ鈋7a�`(�l�1ʬ9 .Oޅ�����AF|)��H�&vl8����'β%�n޿F���'+�C����A�.N�$�fΟWƈ��##�4h�I1J�y""gL$��a�f�`��ࢁb��5CEJ[���G;V�(;pe�D��D)�dQ�g��CזhC ��n�$�>�]>��X�cm�;y�@K�̝Y��C䉈q�Q��!�z-����Z������O�1�Q�6�ɤd@تQcA7�>��<�0�W��P��!0SQ �)��'j[�Y#ѩ
� T�� iF�$ٜ��ff5�d�Y��>A���*���r����T� ��,�S�9)�t�7�p@]{r��cٸ5Fxb$��BU�4g�h������N��?i /U�N���R��W��%(2��p���)�	�o�y�CJ�b��{b�i�<���aZ�X��ؒ��	�G��1����l�����Ý)�!{��)'<ሎ{��M�J����^&��-aX��ȓF�.�s7�J#����'ŏK|4i�۟�pr��sܓa�R9;��	�~�~Z�y�=��g�p�Q��C#<�Rmk&9�O�#�bK)H��ҷD��>�f�+��s����KH�Y��ɫ7葷^��)��ʬ0ź��? �-����'ř9G�Ez���p�'o��2��Ĕ��G�340��O<� I����Kt�Z�mj���KГL�+4恞�a|�$&02E�4�z�|`�,J
�b` '+As�y�#�'fM��ʧF��U�4@X��o�m޴Y�c�zU!�d� f'�e�@��I%������U��c����KŘ=���b�E #E"&��&�3}¢�&��qa�K`�t��]'�p=��}F}{Ӂ�"ؚ%����[Fb�sĖ/�q��[/\�a,V }�@m�V��0w��x�%Czh5:ҍ@9I�.�G,W���'����4���XBe$��L>!��4'�H��ie�-{��r����J�r�q��U�P�1��)�-e��E%��ZqZ��H#o��P�yʟZ�ݫ'�Vi[��
�xF�g)Ѽw (B�ɐ\\1̕s�1
�'�%GbK��%��_*ˎ��'����v�� ��'�,��ǟ�a���Ձ��=+	�C���yR�̴E��at�N 6$|��m@��]���8��bG�.�p>90*�!|s�c�5j<n�S�*XU�'�F�0�g4c�l=�B�׍6�Z�'vǴ\bR���	����5b�I�Bx��d7��q�X�Zi�,�%�� �l0�'�j�����G� ���ɭ����q�`�P	YIb�@DPnq�0"O�5���ۡa`�	���W�Ȧ	�e`Jy8��'?�eB2E�ØϘ'@*���	!J|bM�8�"	�'v�З��L`Jt0�`Q��i�)[=��`� �T'S�����ǍV#�(�&�޷:�4�rh�n%ayRE^�/�Bh���m\�~O�u[w@Y�(���Ô��6!���wվ�I%ʣ5Uq;���,Z1Op9���.lڠHx��	A�'n���֋S�D9�퓖�E�/!�$J�:��]���~'\d@�l�gs�%���u�'�>��� +gN��- .�p�E3pLNd���TR���t���Ф�&"�<�ȓ9�z���,�:qsFx�HˤH$Q��&fd� �$Xj h$�A�J���ȓ�X�S%�ӯU�5lP�}܁�ȓ}xH���k�iɡ�S{�rD�ȓ��HX@@�9JB�qg/�X��ȓ!D������+e�R���=1����ȓz�U���_�"��@��Y�#�b��ȓp�r����h���
2(�I�ȓ��3pG��{�.���ؤsFFфȓy�$�4�wHr��-
G��t�ȓ)��I�@`��t ��Y#�[�6@���z��������0̊>�����+�0�2Q-'���؀���K����ȓ�jx�hŒ%�<���iD7m4���k�0M9���-k���)��H0<�bĄȓ -j @b�έv���*5v�FL��6�H;�k�!~��
D*��Y\��ȓ{��1�1
�{���!�I�3�u�ȓo�.��g0@`�95�C�5V����P(5�C>dѬ���,�
 4��ȓ,֪��ԥ�,)��ӳ��m����$�R�Z��8̄@�"�L�@TхȓL3l5ԭ�u�J��T�Y>"؄��ȓ>��0@�I k�~P1��e*Їȓ
D��������և_�0��s�X��Vs+2\ҍ��(%D��{��H?_Y� ��92q$9D�<���RI�pp�b�ǔX���b�7D�� � �gC=4�JE��L���@A"O���!˗1upE34
?G��}r6"OL-I��яd�<����Ѡot6EH�"O�x���ͪo5�)��]|�{�"O�hn��	yf�H���zA4�'"Otɡd%мO���/��a;���"OL��#nS�s�%B �7h,�V"O4�������3�/�RV	p�"O�-x0��>�̑�MգHbn�aW"O���gN��Q|*ysA���س�"O�� E%�2U��	[@��($�R�@"O&e�u��7a�h0�a�|��[�"O���� -5�!r���?R\R,�"O����g�֙������w"O���#��!�|�覇��]���	�"OJ���%��%�^Hq&�#� 0�#"O����(��d�~QT��NE*g"O��CơW����D�T.|%̩Sp"O��t&މQ��t�Ņ�<ڜ�"Od�*�N��?P�@����9U�<��"O.|hƝ�E6� R�#Y�n��`jq"O�t���/t�bǡ-JԌ@w"Om��b�M�6M�A�Y�B�Ft��"OnВ�ٝJ292���
մ��e"O�Ң]�45�D��I�.{���"O�K�G�o�d|��E 1��"O��8��>���+C!�&!�|,�a"O�� K)/m ]�я�*e>6��"Obe3e]|h�)�߻\�,�t"O�͒�l�w����`X;��ڐ"OnY��p}8�*,́C*��y�"O�(p��8f\���A�D|�"O`X�E&V�7� �9�m��Vx�Z�"OЍ�%P����3lф<>�`"ORii5lM�k��,i�� 5$�^ q�"O>]�s.G��:����>p$� ��"O0q1SX�AY�p���'1���"OĘZ��͒�rYҦ�O���c�"O^x��7��(b�NG�h����3"O�Y� ���B��A���� =�4DzS"OTM9tѨ,��p��
"((8�Ӱ"O�&,W�9��$�4"�Z����C*O�g%ˠm؀���ȨV�x0�'s| ��
�,�f�Ô+A=�`Ĩ�'G�,�q�U5��Je�
�<?����'h�@� �y��zL(G���'C�U&��,Q�9�o!N���'�P(�SfS/<��j%h:ki�i	�'|P|Pw�_79Z]+����xԬ�Q�'��q�����n�HfLO=�N�R�'6��!+�\u�Q��d(����'Sڠ"t�(og|0��ᏼjZyP�'�X����� N�x��G�vT���'� <kv�ܡ:$r���ڊgq�,k�'�p"�^)9��)�"d��(�'7l �S�Jj"�����`n�9h�'g`%�珓o'6]���C�X�Lā�'�z�"��V�J��aP�l��L�|\�
�'`b��G�A�u��!� S�IG�Yx
�'���e,�̬S!"\�@]4`)�'�̡w�J���Y���@��Ti�'�)��ŕk����H�.5f�*�'ъsfg�_�F���]/!t<mB
�'�֑2�eZ�,�L� �	Q,��d�	��� ��9��&��"A�oHr�:p"O��sU��X�PK��B��,P��O����WWN�v"�%4�J��h&:!�D_&8��	<F]Bb��;_�!��#ǶI��H�)�J@H�T�!�D	�Dr9�a��9�-X�g�w!�)S�t	@LB^���ڰ,H!�  ������y���q����E:!���L��`�RO�n�YwNb�!�@�8�z��4�D�R�#�6�!��r_]�w��b�(�a:.�!���;<�6E6`N��08��O�6wX!�D@���Y� ���1�����{W!�d��f���Ð�e���Ƣ7#!�ֆF�00A���@��+@.#!�i���ԯQ�y�r�J!��h!�I
������' j�X�#��$!�D�H�A�ܿ7^e��hՐY!��$��3���H��{u��"2!���a�܅��`���X�I��"O��
�n�>��څ��~���"OD�Ka)�=}�|Cge��L�`�"O��1��P6W�<�sFH�팑��"Oxx���B�����d	*�NX��"O<��r�3�.�0�-I���PQ"O.Qx��w��1{��_(#��3"O�� ���	�\ ��
T }$Ԩ��"On��q��c3x�GJ� X���s�"O0�t��yRUѰ��qK
9� "O�� sK����i���*����"OAkb�D�c��l� %6FU+F"O�Qs Z3N����E$�3����"Ox$�5,I� ���Î4Y#��A"O����'�>Q(pbI�Wh���"O�	Ң�hn;7l���;�"Or]j����z�#�
Ke�h��U"O�ؒ�C�8�X{r*/7���"Olq���8R�x1w�I ��i��"O�L� �����0>x����"O.�+�?k�xa��Dt�`�"O�mIV�A����GmTr`z�"O��5�J�L��i�$�&b�j��"O����-����#�� ��P&"O~PSU��d���U*��(��Trq"O�PcH�3PC`�U3�\��F"Ore�E��&mD]��+��գ3�O���� �zr
q
r��q��}:d��2	�!�D]�u���o����� Q�!��!�.��0eaP�k�W�r�!� 3��p��cIm��W
�!��!�t��.p^f�6�D�\!�dZ�>lz��
�G[�H���
,^�!�d?�&Pi�G��
MV�����v:!�$�6w.A���8������5[%�x��	��9iF�V=J
��P%JFB��/0����Aڂ@yր�P-�o'@B�	�a�M@B��>��M�Fa��n_jB�I�d8J|�nR�Y��2��ɗQa4B�ɶkp1��P�R�����܍(�B�	����R�K�ZX��/�C�IC���`ӧ=�XՊdO�(<tC�I#$�>m�M  �wHD�}�F�$<�S��MK6�V&ˠtPFOϱA8�?D���T�ֲ+"�Z���z�ɹW=D�� <U��$ϔs(�BA�/`D*ѐ'"O��*�gHR�8h2�O2���cC"O����]�i!�@{�� 9O�H}e"O
q!!�B8Hd���ޛ8L�A�"O���`�*E ��h�,�eDL��"O���4�2
�����
	k0����"O�T�cзφ�
 4�次�"O�Y*�F��g"�0D�;�z�p�"O.�I7%S�F@Tt��Mׯs�-�"OZ<�b-:LV�Á-$���d9�S�'#+L�se�X%�U3b@_F����\9H�p`��7�<Г����|Շȓy��s�.��#�8�0��M����.Č�˷�M�	6�U�YR��܄�Ot��WI�O]D�sk��T��'mў"}���4)�i�<T�h��C䉫WI2e9��E4A�� IT�8�(B䉷�$`c�A�&����g�Qa��C�	*->���eP�<Ԙ�N�t��C䉎y��Az��^�y��1͔��C�I>����D57B����	bn�C��Y�$�
���)�L�`❌��B�I��<��g͎@�Y�&[5R��B�I
B�<�j�n��1�g!�"EL�B�		,v �rB z�<��ŋ��)X!��!�b���ś4u���E2}!��Z����߈+*`P�MQ(h!�d��:K4.� @����-�+5V!��
���С��4z9L}q�VA!�I2
K�B��C-���‽%�!�D�'�ݢ��L/'��{�$�:'!��M?�Z����+� �E��^#!���j`�u�[<1$E�!�DE1�L�Q"g��W�T
ă@�!��	|x���ĩ��!��`����F�!�ѯ�� �+�%r�J�#�,��h!�$�O�2�ѝ7Yy%��(�!򤔙DT0�a�֕|�|H8H�!�dX�V���G�T�=S�ѤF�c!�$��B���G��:}�5fʋ)!�d#Dy.�q���1��p��$�!򤐡6ލ�� �G�j�c6��O�!�$	�nܸ�����QвT���	;�!�D5E�v�I���8�а F_<�!�$�V�`"�Q��Ar�2�!��AN�lI��D2 ��xK�hT��!��
�mzDjb��1~�y*���!� N;~�`�N�'�6�yF�V�:�!�D�5O�ܔs�C�<��㣓�-��Z�)�N��I�9vJlx4�<�y�) ��D	 D� lи<p���y��F0쭁�kŒ[/�0(�y�%]�%u��H���C�.4r��L*�y�G�^
�}��R%,�1S�lF��ybW�j尤�
y�0q���݁�y����N�feY0l��j��i)1����y���A�AH�aOi��"a�H��ybX�y��#kP�g��Y+ �ʹ�y�n'||9SFȂY���(� �y��\����n�L���)�ʔ�y�+��R�@y��Á&3H����똞�y��F��J��̢#�i��y�#�>m��9
fR�#E�y����yb��	 +ʩ���&�61[7.ʺ�y
� ���2�2.JT�gAU?Z�\�;4"O�-���+%B���B���}�;�"O��� k���a�gk1Gz�u"OV���(�1'�8�4iLE�4�p"O��
�pKp���M^d���"O�]��k�D� �-P48l5��"O�Qcv�D1֚���Mا-&�ɦ"O�iۓj8x�u����R���{p"O�heă�?a<�H�o�i�&H�O�<y��%��������/8"�n�L�<)��ԀJ��UB��M�!gcMI�<�0���/�<��&�FP������LB�<ِH�!z<4��aܜDt|�p�D�~�<q0��/whɂq�ݱNV(���}�<aV��$Ϙh�aOi�=rph�|�<�O�y�Ta�@,�pm�'�m�<1�ǧY\Hy��S �$��7'@b�<q��C�Z�@dr�i�#z�}�E�v�<9�L�𨼺�ۇ+"d̒B��n�<agQ�����L��/d,	:U�Q�<��/U���	iк��	K�<�G�O�rԣ!M8:z~���I�<i�@�f��S'��M�:m�g�P�<�blƢI�r���M���"�o�H�<閮T� ��eh�nӜ��yZu�E�<Y����"��WA̒X8R�K�B�<鶫�i<Н����6H��e�]@�<!g�u�����.�3�&�y$F�{�<D/vZ��EKJ�o>ڰy3ϝw�<)!ǆ�6-� (�@��$��$)�lK�<��o�7��u�T!$���b|�<�c���P�hqq�K�w�f�(��OO�<�1,
�2@
���+�EW.e�֠�P�<yc��5#ݒ�Pg�)e0 ���H�<yQ�ک�d����S��3G�Do�<��Ԯ
0��m��l����ժ"O�(�S(�X�$����0N�u�"Or�"��F�:��9�g�AF&��"O���L� ���$�ߌ;⼱�"O~P9C�%-`@�z�Cʾ{p�u�6"O����*�'49�(����;m��B&"O��s���S�����|�|bc"O���g�;hW�R��Ѡ\b��"O,Q3O�a�,Щ&ύ�ZF���"O�H�'�ԑ?�"-;�(��g?v�z�"O����
�%q���(Iׄ\�ƄJS"O<)"���z)ܱ蒪P^���[$"O9���*l�:�h��#�����"O^a��:��y�B�E7��(��"O�Y��ףs�]�!�ǰ6����G"O�]I�
H,.�6y�ƈ��xD�*�"O�PQ����Q����t�L�7"O$��h^�^�`�G�H���*"O� k���!��UЀ��f�d���"Olq�铪'�����+��f�&��"O`�����e��I�� C�^�j"O¸j�cC�5p�2��A
}i��'"O�p�V�#��a�Uk%IcF�X5"O��bq'A9��t"��wM�y��"O�H�Aӎ)�:��WF�*w1~�"O���G,0���)��kk=P1AB"O������$@+�-0���"O�����Q�l��zP�Gx��a��"OVK4OG/[���� 荵u� ��Q"O� ,X!�ID3{Mh� ��I	]���4"O����Q
u��5Î32,I�e"O���6��ZR"��c�I�L���"OPY�*J7]��	��A���p)u"OR�qsDʠV�*��3�O��~�	"O`H`#L,g�Z0� �-G� D"O��KЯ4"�$�Y4��#2�٠�"O�� pK�����QS�C!E�9
!"O T��
Җ!�x��2�M(ժ���"OX�	��3�"�i��Y$����G"ONp��	�([F`iۚ5s�<�8w"OuB0 ��1. q8��9��؛"O�A`�
�?�Bģ b0^�@"Ova�T�@��J3bgS%9��2g"O6q�ІXIT����Y�|�L�y�"O&@��!��3���C�EN�^�N|��"OP`pud���~��'d�'5��"OfL#��U� �]q�Q?n��a"O4�A��=;&�@h^��\Y3P"O�U"��U#l[��	R�˿w�T�S"Oj�g�IXZ�K
�n1��"OƁ�D���(;j\BCə/�Щ�"O�� ���n�p�khq[f"O.!���9Rt) �M�ye~\;B"Ol�HTlR�~@�p��]1#Z���Q"O�dD��i�l�[�-�5%FZ��"O��S�b�"��bL�H�4�:�"OH�eW4�A���cք��"O4,����&�����V�kt��(�"Oh�BQ�W�n>X1q/�]�X� "OL�P�D�>��I��gƔp:�"O�q&%ϗ.�(�a�W`��i2"O^����(��Y�7B]!r/Ҡ�"OH�K��:X{�!�� ?&.��"O�aE�4}R)�M+	&��f"OhI9�eW5'k��r�.R���Q"O���fh�/���s/жp�U��"O��H%��!���,TW}��"O�i��
W&mt�,�t�A�ᓲ"O&< �M��-��aY�K�x�E"O�K�)J�6��,�s�����x�"ON��`��c���`��.�^�K�"OX9��X'rH�ت�/��8�l�P�"O�E�F�th2mc ��d�X��"O��Ɖ�*�R9 �m�?2z`qK�"O�`��:)I�	scb�k,� �"O$��Vy�@�6�>qOJ��"O ��`e�\n���b��j ��"O�����p�(���\Z�[p"O�E�t�Y��D�˥�A�~H���q"Ox�� �mTe����:��za"O"���^�y��-��e#�Y��"O}��IT/J�\�Ū��j��u��"O��P�+���OV�-7��v"O��"�^�an���O=+6���v"O�Y0��K,� U������*r"O���r�S�"=T�;��I5Hhdar�"O��`g劵K�M1V*�W��"OXp��
�)@��V�˹l_��"OI�"D� Wc��P���	Wy��c4"O� � '.Xn�0[S�!P_2uC�"O�5��Ș')�9QeeÝ(n�c�"OFqs�$
$#����1
W�S���y"O�p�0b�E9>�PX8B�l�t"O� ĽI�ZQ���z0fK�%(���p"O�E
U	��%��`
��C	}'���"OX-� �	�b� S�M6 ��e�"O�U��XQRē���x���9�"ODr�Iދ�bbF"���"OV��hR�_�M��V�]^��"��'�B��;�'oL@���Z�(�H��!/��Y:�'>��Y��ɕ'�"d�� ؾ,B2\
�'��!#�N�hP)a�'H�(�	�'a `R�	�&_��R�ւ	 �3
�'��\�f�.W)���E�G2�P9�	ߓ��'�Y
�р��FD�(dT@	�'[�d�r/�-[��3�ϩ-,�d;
�'1��C"5H5�x��ػ!x8c	�'n*�a$�]�;������%�	�'�Ұ���S��!Ң 8!�j`��'
eJdH�/r}�ɚ��Ͱt"O�U8��ʇ���yw��#ڀ��'�b� &�h`�t�@�k@��X8�!�C�7?��� KM�z"�uB�@>N�!�D�J|R���0B�f�
a��n�!���7���C%H��qQl0�!��� Lʨ˓�Z�M8 ȒC*0C�!�Gh�x��6+Ft�7 	i�!��
�/��0�c��RޤHZ�`�,l��{��'�I��@E!��Ъ4mnX��KR��İ<�n�~�C�%A=w�:q�Өȵu<� ��`1^L�1� �C�(|ٴ"�3ikr��ȓ?�f�K��K<v&�@P	�2oh���ȓA��7��W����q��D̎$��it0|Ir��B�	�������)�ȓ;")b���:�t�Xr�Fn�)��	j�'d���QK�����׹�������hO?��̃L��Q����Ra�V��H�<�c��i5bI�Ѥ�(cu6=AiD�<�	ߣP8��Y�/��fv=bƜA�<A"��s��!��		|�
7*]~�<�P%�T��1�%�>�zf�Uq�<��,����1���pR�3D�A�<2��'��p���B�I� ��L�'��'��Of1O~��t�_-���	�!��[�p9Ȁ"O&P�/αA��,Q��� 9��M�2�'�ў"~��o�Y��!�D�W�{� ��6����5�O�I�żq̊*!\�@�F4�4"Od�OĮyIĀR嚹�"OVl1P ;F�.|ʆř:����"Oz��Х��h�� ��h ��S"O��Q�)�2�t1�d�	)Vb�[v�|2�'��e��ン*�2qK&l��,�����'� ��C�,��C'CK�
3���Є��K�ư����[�zx7J	�qp��ȓ*� �燅rD�1����hj���Zv�	W.*HV�z�}�\݇�Of,��Ò7Wu��ʲ�P�%^���j�B@��؊���b�@%��ȓ9�DR�D\��v'ڒe{pq�ȓxe8��C�Y�^�̨
�&Z�"� ��ȓJ�����F�	�4�w%%Vd�����&�I�$֤"����7��:Ų�ȓb�%��#0~-��m�.L� �ȓy�T���	����ju�J�8V�ȅ�IX�'^�lJ�&ئ3�^��E��N��EK
�'�f��N����Q�Y����'�F:p�	R��%��fL6T&"���?��S�? \����O�H2����,����6"O^�Ҭ�>�00��n|� В�"O���0CJ�3�޸�c�[�4^��i6*O~���O@�S)2A���-��d��Ir�O�LԨ �V�Y��e[''l��'�� �6��!U4D��T��zZ�j�2�)���(ot\�S R2G��ͳqb����D�<�
ӓ:L����T<v��@��؄)�Lч�GK�L;�LN�a��C�#�	<�(��&s�B3��B�T8ׁ�.a�d��ȓq�(�����0b�8p&��A�蠄�	�'o:MseN�C@���A+"���'�B�Ѕ�@:�Q��,B+=�,lr���"��8�!]�����
EbXd��""O*]�av��90#��VJ�@��"O�� ��τic���W�VPdj��"O��� �G�J̎���]4� 7"Od��dʤ~�����
[ �j�"O�LY�N�2
Ā�E�eA�)у"O��`ʊ�J��d��F֕91(M�F��wyR󉛓W3^	��ët��@��H�:2|!�]++���\Y`���hޞ*��ȓl��D�в1�Υ��)�0ypn��ȓXY��0A�	�??:U�s)3�P�ȓ�:����év�
����Ox�X�ȓc�P�2Qa�0'j=�o��ԇ�Y�L��.�k�V�k���{b����p6��'�x4h���t�v��U<��C_�mkP<�ƌ��t#����Dl�<�so�:&��s%�N�̤���B�<1�L."�x�� SU�d��ʙA�<��i\�Vl5(�lr>x���y�<�F�Y� �4�"�����se�`�<QA��8l'~�#+3�r�C�+`�<��bʨK��LJ���T�S�]]�<i��/F|�t�u�ڦU�@�6��[�<��s�E�2*�P�p�LD`!�L+2*]�D�^��8�Ь	�VI!�Eڶ�Ju��|��Y���I%N!��Yu�����<s��)Q$G�C!��Nw���U	O:ncj�K���x!�P�u��yk���:8W�QH�Z/1P!�D�)~;xL[���)JN��:�C͒J!�$�>r��&[�^LZ5�X�\!�$����|�  ���%	cR�,I!�X��L��Vw@h�S&S�!��M�&��'�C�T�6��m��!���x�N�xJ˂X�qb���'��Q҂��7����/�k(R��
�'�Q�4ѢB$81K���3���
�'�l�nU����YfL�Z��x�';P�&�s���c�!U�,Y�'�J�i�LP���!N8M����'��\��]��2Myo҅ ����U��F{��9p�rȹ&��~�~����Z�
C!�6ue�TR�ƈv�`8qP��<S\!�_i�ۧEí]�x �OGI�!��շ+W� u◈E�ޑsu.S� �!�dOT�����tduР,P�6�џ G�D Y�G*����<'����� �yҪ@(El���÷M"��F#���?i��?������"w�X�`r��Sg`�H���1,����0)��i1~�n��e��
�ȓ t6ْ�m�>�̑˥��Ań�S�? �ɸ���A�CѣO�R���"O����ڗ9U���爒#��=)����<ُ��ߟ5V��a��6dN��H�!�䞃E�hX��L�-W�@t( ��b	�'����	E"�8M �4� �YHajR"O:@�Q�D���
̲z�$"�"O,	9c���c0�0e��C�z�h$*O���*A�E�z6��R+���'(��S.(2�õjѶP \mK>�������O8���a�.w��Y�`区K� ��'�Z�!�@̯PT���2�<vmAL>�������O�@
1��Ң��!S
��
�'�H��4�̂#��,sA,�+Pπe"
�'���q �a]T5�3���Dg츊�'��	p1kׂv��	r��=ZtQ	�'��m�!	ԉ�� �/�@�pjH>I������O)�)c�
�a�2���ՠ>�M/O|�O2�}��?��3
���2�.^"<)&��G{��de�x�Dp�E�YzH��ӎ<�y���S_��2C�',���+�y�B�ծ� .�;)\��rR��y"���h.
��Q޵'TP��1n�y2ă�& %C�`�9%wR�@1�P���'ў�O�0�H�l�>ouh�Y�6l�����hO?���/�\%���)pkRH�-
p�<A3m˾0?��x�˝�<z���uITA�<�@M4�Yh��
�Z�桃��c�<���Y��Z������ LK�H�a�<!�[�$�����F�Bg.@T�F�<�F����AIelV<mT:��G�E�<Y�+юc��E�1�]5u~T�r5�@�<9`�S4U���J��X3��`�����<�Ӊi�4p ެd�d������y�H�E�I�.��_�����B��y� ,0x�� HϣF�" ��-�y��ۚ%�V�:7�CD��i+2`�:�yBA^�e����� �Iz|XAlֱ�hOp�$�OX#|:�U����c��^%:�"��[�<�6m
�=�f��&�7`a���JXt�<!�*�8���b7W?N ����U�<��"u�����kK�+ �a%FLT�<ن�J)>J�+Ɖf8p�̄d�<��A�Z�\�/�9qԅI"��k�<�C�
(jT�!g\b�0d�'82�'#1��a �{�$������X��"OL���cS�t�v9�d�6~88C"Oΐ���:�������1��h�"O(�3�d�5b����Q.R�r"O��Æ,@ xr�8S��cM��U"Od����oVC��)u����"O�������+V��Bb_6h}l����˟��IP�O*���Ml�pnU�j�9J�''t	+G��L�6��	6Cl��'G�l(���'<:N	9c(_9�`��'W�웖H�aR	"��G0c� ��'Cf��U�_�G��;BcN�(�����'n���"�	�2E:4��nT-i���@
�'�N�yp(Á1Bશ��2[g6�Z	�'�>U�c�aP�x����+(��a��'�&A��b��|�es����&b�����d O
5"��#�4��M�&!:*���"ONpyE�&$FP��KL�x@i�"O`5h� �g���;4�S>g&�pZ�"Oƕ[��< �z���.��T�"O� ��v���~LU��*L�
�^���"O1f��m?�]I�� q�$��vX��D{��	R&C�!�3)����H�±A�!��';Ҏ��6�ޣ1(�]�4��)p�!��W"`$���gD��&e�j�S%!��^p#�)� !�g8���Ye!�Dӗ<A�F$4G��� (߷[!��<�b]kĮĖK�L�F!�d�	w�٢��	��V�Yc#�5#9!��Mg^�꣣�Z�$�!�3r�!�$�*�P���\)K�ΤA_�!�$� %T~� k�1�P��Ģ���!��׋ly*�B��AZ���`�-Y�!�D����U�朤KL����'c!�P�.�������:X�(�u�VQ!��rl˵ ө
Vh�2*K55ў�D{B4Od���/�=V����T�Ȕ_�D�cu�|r�)���Z�F��.G��R'N�JFFC����� �@�g4��D�R0C�I!5���2�N`En�"@KM�B��6�f!IVON�"�F<{�hK+ްB�(G4�2P,�)C�����u0�?)��I*@��(!AL����
r�Vp��D<\�T��^;E�-�qIO-ԀC��/E�p��#+2�]��"O6�ZY(ԉ�^,*��xg��T�!��U��+��Eh���Ͽ`�!�Ny��4�C�V�a�4FT$�!��[5 ,�z��ȿvϾ��teK�Qў܄��"`�:p�gK�A�iS6A�*�6C�I~U
h��V�GSV� ���%VwC�I��攫���0�����GX1�؅�IT��i6\T�ƂU⨕���1Ҷ"�5�2e:4�V�4�����$:�	��f�)B�X�I�b�����囂�)�lY�k&T��{~�IA�������
� }�Ɠ;!��.D�]�~)���T,��di��?�tBk�\� ��.yN�� ;�y"��9^�����	z`@g�ҥ�ybI�zv�T��rf0��q�0�yR��' �6)�7�Nff����J
�y��b1�@��eZdn�\�f���y�M�>Dޡ�2�T\>��䤈�yʖ6E�%����P�e���y���;�\�A��Uw������y��U��<G�:^�]��k	�y��D�}�%J��1u� r�Μ�y������P'b�����j_��yb�P�@��)�(�E���(� �yRDY�E�ؚ%�ػ'�m`嫑��y�眑f{��
x�԰:�A���d,�S�O�fY���ĺ�F��%��C����'�Z<p����m>�i�(� @d1qH>Q��?9Ói�����oM�*2���%F���,��?N�ݘ".�vª���*b�^��ȓ.wjuc��6.���y��Ӎx�JĆ�L����˲O��9Z�A~7���1���J�ɉ�i��L�a'Ʌ>�&0�ȓZ:�JE�6xF� �V�syL��d�&H1ć�8QZp`D6�J�'�x�'rax�TgoV8�����a�S�O�yB��7�j��G"��y㞭��+ā�yb��v�R��h f�b-)� @��y
� ��b�ĭ(��X9Q,F�+þP"O4�G�'�h�rʌ�2n��"O��*�,^����1 �0y�<Z�"Ol�q#�7���x3��)^�`���|��'w�'��X�ۍgL�b@��;(��*�':0iY�nC�b���BeB8o����'�Q�%�O��M���1�]a�'�� : �=��9�`�;z<|yQ
�'�ظyUF$h����5k��3�'�����l��*�2|���K�a�H	�'or1��G��J]�A0c��p�<�)�'^x��$��}h�YW�քf�� �'+��h�V'߄ɧ&���(��'����e�:7��ibd�1h�(�'���X��"nR�I�a���ۺգ
�'V��U̝\��}�`ІB�
1
�'�T#��X8��jA->>n��'�la�cl�:����e."�J �	�'��b+�
��Q�7�#����'p�P5F�*a�u�ƍ�4(:�B�'�4,R"Z�5~��ևX-�t}��'�L�[W�մ٨y�p�C�
�m�	�'�L���՛HH��Q�� ���''d�����GZ	@F��{�v���'H$Q` �A w8�صA[�E����'u6�� ��Dڀ���>;y����'���8�"��S� �4�Y�1���'��pʠfQ�Uy�a���=!z9��'k�R7��8M`�@������[�'���q0ώ O��	��(��E~Ţ����0=1g˾b��d���?�3@ �b�<�&��,�"�Qr��(($�d���a�<���&^&0�S#S#_�(���B�y�<���C�q0�EK�}ƌ�V'�v�<1�%8Cm���?
~d��rj\~�<�SbǠ,��D��:3ڨ �q��w�<��ŕ>�H��]|�>�r@��[�<Q��E<jFՋ``�%uD�����V�<���Z�M��)f�]��)D���5'�{Cj�B�KI�gm\|��E)D���q�M�S�J��Q��!J�2ؓ��(D�j��	�a������|w:��so9D��0c�Ɗlb�tC�@�2!�Lx8D���ck	 F>L1H���8���5D����e؛z),�rq왱$fn�J I3D�TC�c�.C^Q閰8�@xj�5D�d�3"6�"@��G5 �;&*)D���D��rh�1�gڒ�:��$(D�s��|����2O0/� �h�(D�xU���7A^�#E�� s!��:�$D��1�(V@бBu�Ȧ$������$D���Dɘ>`��2�$fb��m!D�P��ݝ:vUI#+ؒHE��H�"5D�<���C?0�~�Y���#!�4i�g.D���$K�M�B  �+��S��\k�/D� )�)A�ޡs�D�
茛�f,D�h!�"��vH�K�`��,M �E/D���EHF(c/*5#�mhX ��A.-D��3��Z�N��Irn�4.���*D��QI� {�`Z��j�yh4�4D�Z��=d�Ɯ*���.X��P57D�H��T�Vvft��Wn��e2/4D�dE�����,s��V6 ��d��b0��2�SܧE��A�H�8���ℛde��S�? �\Z�勯-�$<��Ǆ�DJ��j�"OT8!�nE�Z��9s!��uJ��;�"O)�AkGn���Ե'1��"O��K�m�=V��2��ɵ\K&�� "O�q��©VB���E�K�b"O^ic���7U�b�%W��2r�$)<O�	P#b�7j��(ࠋd@|���8D� �D3;�V�)b@](=�4X�3D�T���Y�a6��Puj�p���AE6D� �&C�4Z���Z�%�@x���0D�|r7�צg�()��Q�~`�QI-D��ӑ�ſY2�\8h��M3\̻aD+D��� @	�!nJI�6��2.��G�O"⟀D��'��$���QN�X�2�F@��`�d7��Zr&�(���:'
�gݢ��G%D�Xv��h�6 	1-Q�WFH��"#D��R�`�\��y���x
���=D�,  &�.6.�"�!=���S!<D�\�Dh�G ��x���l}6��:D�`Sq�a�~Tsiɾ��Ykc-�O��	�nu[���8bc�c&��7VP�C�	9hg�])�(2'cC�7�x=��'��I��o��fmd]��a�4;+.�	�'_���@�H�2Qڍ���^|��'�v��s��~R�I��kWA����'�\����8{�)��Z�'�qK���0]�X���T�F�����@%BT�ƪ;%|P����S!���=DHS拀=  �q��Q7�!�$� &OH�ƄY�W8��w��k�!�Y�[X����U�"!ȕ��[�!�$��L����%��V��ReĔ�!��ZLԀJ�)�c��]�t�M|�!�$��f	;��	7?'��{p- �m��ID��ΓkId@��ɇ/���HW�V)v֍F{"�O!ֱ3�GH�?l@�B��Fu*�'�
M���[�mԠ���֚qeԈ�'i ��� �ld@�V�I�'n��$�ā��:E ��;��;�'�PͰ�%� ���̲/m�h�'��\yB��*x��Т&�f �,O��D(�O�8��j�.[2q��K�M���e"O�dr�/
�^��:�<��'"O �x&N8�A��U�%�$��"O�H��Ň�]B�J�CĨf�(�Kw"O�l��N�#��̆}��
P!b�<Ѣ�v�D�ׄ��r�$*&�u�<�S�J[���B�4i�ʱa���q�<ɓfF�(t`�.�1���'�Byr�'OҐ|����
Nj4HZd7�:-*�e�N&!��مw�X8�b�4w�V�%G�
 !�Dܓ)��й���8?P�u�pC��b!��56t�6�R!�)�� .O!�Du�j1�%��1m��l[��
�'(�X;�j/$�@4�'��c:2m��'��9"�F̏3j�4�E�/W-P}���hO?K�,ք�2� 3�U�ZL�B�RQ�<��Ď�p��d@�
޼�b��C�<����.m�ƽ��.��jr���dB|�<�6��E��E��ɐ�O��B�Py�<q��@�c�k��\P��Q��q�<�e�Y&S|j|�p�C(}��ل	Uj�<Ie$��H��4b�D$� �X!�h�<Aц��R�!��\@B.�]�<� ưy!�ۍ �8Ţ�C�6�ȳ�"O�%G��cn�iHf�9�,��C"OD������q2��㠉�oe�`cP"O��&�U48���0��.HU֩�"O���L��*�½�g�� L~q�"O���!$��!�θI�a��H; !"O�	�p��:N!�*)Ԛ�f"O������hf�8�d���k�j|��"O��MV(*�B���gG�h�����"O�E��hW/U.�ru���~�u�"O���5!C>B0��@V�6&phE�"O�|����4tб��$;Qe��˲"O�5��[2�L��)&eT�-�6�|��)�ӷkb>xS�bu*}aw�-Q�B�	1_l���'Ǭ7���r���)j,C�	4i�]���'$j�p1�㕌Ew�B�ɦ"���pfiP����d��Y�dB�ɲ 2ȡ�)�S �E�e�PT�C��9v-�D�� �Â��0��"O�Ys%/�)sL�R�X^z�����'�S�)ĿɬeyŴ�=v�Ii��
$�!��Fc����N� n\9���ķ^�!�+Eш�C� 5Mʐ`�%��lP!��,��A��e]���<��Ӄ�!�2{��
!��������+�!��׃� ��]#E����X
�!�,Ӵ���gbOƌ�"�ޱ;y�O��=��Q��eE�[+D#�Â�*��Y�"OR����+݆@��G�(��D�"O��	���2D	����1���F"O��)0�4{T��0o�:X�@9�"O�`�5 Cn ΜC�-��>�2��"OBI�a�W^�N��n���"OP��b!N  ��*v}-X8!0"O� q�!J
� rl����D��"O�B�"G�2?�Hc� ��)���R�"O 5)*X2 �)`�`��7"Oѫ&��g���Qq`�DR}G"O,����2~��хΙ`�Z���"O���&]�G�D�e�C)-���#C"O���E�I^��W�֫7�.�5"OL��M�-=���Ye#���Ĕh�<!��ͯ)�8�i���j�أ�EI�<�������0�#���s�=I��I�<��&�!j�=ɂ`8K�|�r�]F�<��i
��e�э[�1P�k�FC�<���úY�ɶ�̾Q��s"΂��TF{��i�wa�\���Ȓ$���۞]W�ʓ�hOQ>�i���5{� ;�끷*�eY�i*D����1,�h� ���$�� �#D��3�	E9RY�d��B�br�#D��Q )-y`�{�m�>b��Rǫ#D�Xa�M�i�N��B.V?�0ᣄ�6D�HQ�I�d��T��֋=���%�5�O��v��	U�
4��੖b��1ƶ��ȓ֎��&�|3v�G�+Z��ȓ1����u�N5%��A2�O"h��؇�/Iܼ(����ekH�6aD5|����ȓg���9���9UR�����r��q��t�V�S�Kt=Q��U�sJ8��"݊�J	�'��I�K^w+й��II̓W[���
$*xA�K�?7�Ć��ه��5>��0�n,���ȓَ�Z�j[9I���������S�? <�X�⁤<���&�A6$�vukC"O�|BD�%3�F�"F ��'� <�V"O>`�B�&�A!��%N�>�z�"O:Q�%�R�`�e�H@����K�'��ɺY花I�$�q@6�( �T%M-�B�	�=q�pREH�8: E��o�X�C�< j�a����*f��c
Ё2+�C��Dt�}�H��HՂ2gɺt`^B�ɭ�)B�b�	�YA�[5��B�	�L�2 ��K�5z�z���C'B��C�IV��	�DQh�W�V�M�C�	BԒъՠ�^�,H�`(��4bC�I!v4� �/�9Mk�%Ó��^|JC�?`Sx#֫T�n����NKrB�7�� 6hJ��x P#m�	:�2B䉝U�RӦ��
�>@�
^���C�	P~,���	H����0��]�C�	x

d!Do�4E���ܶ9���F{J?)V(�'�J<�O=V��+�5D���aJЌs�\���� �l���-!D��@������i#hG�P�~�a��1D��XGF#D�\�
���:�4��e-0D�\�f℺=�1�iϬJ&q�V,D�ܒ�G�O�Q	��Y	A>��9��)D�`�c+��^ N���0P����� (ړ�0|��G(O/��@�D�?g�.<3���t�<Q�HV7M+�u"Q"B�Sx0��A�v�<1�f&o"|�bH��S�^\�n�q�<Y�bɾW�3�" �gc�(*��m�<�6@	z���3����'xP��6�_�<Q@�ȥݒ�1䉆��� �`�<�s�q,0U�w��a�ܰRf+
Y�<��I;5d=���J�
�1v@�T�<!J=�"�!�J`n��Y���T�<AR�U��P:�o�`����$g�I�<��Ɂ/m��+�ƈw}����H�<��߷m4V�B��C r� ���\�<Y�Ӗ���RV|���4�U�<у�K	w^9Y5�߂g���I�$�\�<��H�ߴ���̙8g�l�b^\�<W˙&N3�H�*õ1���a��a�<�"��d�F�� -}��,	Р�]�<��Ϝ�u�N��5����nɀ��`�<!+�T�(]@"m�:*E�lȥcPZ�<�2H�(M�L�[���;9����.\p�<ѐ�_�h3N��r�=w�j��"HV�<����a!
�e�@5}�<���P�<I��.}�
�!vo��Q,�/�J�<jVkt����8
D�H��a�<��@Й9��U#�ė�	��DXt�<a�I�(c�2���ɺ���[āKt�<��f+gܖH��k�,� ����Dq�<)T�L(E0��U
<x���i�<yF�	?Z��P��KT�^_~��u�e�<��l,8�����a�S�B� �(�|�<'3�J]����|�uHCy�<���S�&�BI�Q⋒t�Ҝ���w�<���yÞM���Ж	ވ�Q�nRZ�<ѕE�}����a(��pnP�5PS�<a.;6��R"�V�7�j��P'E�<"E��+F��#�B��%h�M B���$�앧�����1�\�F8���cKJB�I�7.�,(�̈́�4 `�j��=. B�IaKf4����7-|f�S�,W�VB�)� �P��T�P�	�S�*kd"OD��2�	6 2�H��Qp��yG"O�1�6Ŗi��	*w��46�u"O.��REOcp��C�^:{,*!��[�%�PG��'�`Tch-jN�<���F�i��'���B�A?\�l�X�
����'\p���J�^���`N�y	 ���'}�K
Y� ,�-k�G׮r?���'\Bd1Sɝ)1W@���O�"_�L���'A�@P�+�"|T8�Y�Aen���'>l������<���O8gI��+�'�8�0���eDf���X�ڍ�'��� �	t��qg�ŽI����	�'�S+��SN����E6=��	�'[��ha	ϛ_�\D9�׏2���A	�'�:��LC5�Pԣb�>2,�Y�'��ac!��L���)���ě�'/:�8��і,<"=����Eڨ�'���!�]V�r��iW�p`\�I�'<�(��*n.LICE�h�F4P�'�N���"�v�,��"���#�'�dŸ")C�4�5����T)�
�'\���^Sd��#� ^�Q.,�	�'b0"f#�9t��}b��ݷT��J�'���C���D~��"!/�R#���'��N�s���q@�^�H�4d��'���W��5'�<��@ɄBzp�(�'ƀ���	�~��PH24d�Q��'���+ �v&�iۗgF{D�\��'��!���e��*�Ν����A6�9D�Њ�	[:S~V0��Q}�j��`"D�d�ЬR�k�����B%�,Ycj?D��á�U.\٦��?E*a*�%>D�������v�"�I`��2�D��P�=D�p��ƚ�p'L}[�A;	�wo<D����ƕ�nT���p�֋V��P��:D��1w-S�L�PM��'U�+�&�	5�6D�L�s�A
s���[�,AՂ��@/TC�I
p87jQ�%��&��G|LC��.:JXe�e��)��D�/c��C�	�J@(�����z��!:�g�� C�	�-D�E��	8W��<NB�	�]��|X�cԜa��q���%��C䉐_��B��3�dI��f�R��C�	�*`88�)ѫuT��І]=U|C�)V�% �"�� DH��M=u�rC䉧	�Fx�Ūü^�*e��M�1.B�ɓv��C\5��q�CJI�|��C�	�Ҽ�a���4Dp)s��*4�C�I�_\�`��+����ȁ2s%��Q�"O���Q�Zh5�U�xX7"O�i�ÆM?q&��3уǶZ��ڡ"O�dA; e
���̋S@�b"O|Q�ʍj6h���W�6=Xi�4"O��K�se��$��
p&��h7"O���͂*+���d`0"OB�Q��œB�؀H/M7Tx` "OJ�9�,R]nL[�F��X��r"O2����~��1����Lsp"O.�Eł�h)�X��E��p��"O���G��,�"D�I�N�|h��"O�@rr���l���B�p���kS"OH�K���\�:�ᑅr�2��S"O𔒡���,n4����ɒ��8I`"O� �u��DV.�0ې��I��3�"O�!��D�o�=�B鉀F�(���"O.��!���E�@1��E8qr�mD"OFxi!#b���F	);�@	�"O�-�R�V�58�]:�h��,%*1 "OhM��ۨ��yR�ӥ,H1�"O�9r`*<�j�!Pl��i����&"O���@�ӦaN!�2�=S{:�"O��c�M�[�� ��Ԍ*i<��e"O�Q�[�P�P��V��$8�5��"OaA'ʵH�"Ԓ%
ؾB*�eQw"O�ɶ�ME�x�4�"O�l8��G�Vrv9��HW�4)P��"O��B!Y1G��epS.Y4N���"O$�� �]�g��IćȮ? �`d"O΄:b R|�	 � +2�Y��"O�M�篞�i@ǡ��l�s"O�`��1�(qygB�c��#�"OB�{�,��:�#�Q� 6>��"OX�b/��]x����J4�E"O��ɇ-p��ի�d[�w��P��"O.���K�W�*�j�5w�<@��"OИC�C-��|B�*�"(>A��"OH9c��$��L8�V��0�"O]pmF!eۄ��bg�<i�"OL�b$�hcn%��@AK���"O�HÔ������N��\�ȉ7"O�@��%�0Oc�t��-
:�(��"O�i1$�ͽEIz��s�M�p0�yG"O�m2$��K��5������H�"O��P����t_]�f @�Mg����"Oj�ᢥ��T�T8B�r��U��"O4�g냥�\t�]J����	�?�y��O#iM>�w��?��AG%�yr�0P�|�	Æ� �����J��yҢS�c��i��'#8A�$,¸�y�b���2K/zM:�	3����y�HϾ<kttg�o�l�2GW��y�`K5MN�c�S�m�XM�2�D��yBć��$���*k��I�1%*�y�BE��1Sdh^�i��<��ǘ(�yR��+�����n�z�)��Q*�y��t"��5)�8`$ � @��'�y�$U&���kčoS��x�.&�y��3to<�%k
}�f��&� ��y"dΡfw�85ՑoX
��@��y2�I;Y��u�T�ίmOJTI5�Y�y�W�΂�jdj��:�J�a$��'�yb�(Cv=A�(�7����(^�y�d�a�p���Ղ6(j��BgZ��y����C@�f�M�Yf��2�M��y2->H$FZ֨�PA��{���8�yR,U�n�x���:}�@��yb��!{�	�J8�$�֖�y� �U��
u�ܽ3� e(����y2�

l��r�W
'�ư[h���y�Dڗ"�`ɡS��$��H��.�yB�����؀a�ˊh��A�Y��y�B�-l����`�er�*��yr��BЦ��d���b���"R!�y�ÌX^�r�f�*B�োX2�Py�ؼt��V�X?��m��@RN�<��Ɍ(�f��2���\�����I�<��*ԎN�d,:HD�C��pe�IG�<� ��C3I.�(I%�	
b̉"O|K��Ƽ�IQ�b�{�Ѳ�"O��AS͈�wG����K���`L"OƘJf��u�#F�^`<	�V����y2�ҽ�ՉP@O
IhX���n��y�/қVΜ�qEםE�at����yr,�>�K�@YPic�K=�y"&�,��;�$,=��|C �,�y�,��} ����ـ
���("���yҏ�1I�mc�	�Є�4&[��y��"��0G@l�ȣ�L��yb��.t�U�q&��k&���B,�ybC�|�D�7l�9T�(6��y�mOO�� 6�͠6b���ن�y�\�8���[`��3� �����y2�ƕP+��q��w\��fK��y�� (R킂�,f��Q��
�yr��b�c�]1d36�B6���y�":	~:�2ǮϷK�����)�y��!w݌Q�d@SH�hș�����y�Lĳ|$ͳ�	I�Uz�4�E���y�Rca������9�8E�E��yb�C0di��	�d1)qj=����yb%A�A��h*lˇ$l�4�G��y�(�)}�֐����'�����+�y"K�.M;�=�*I�l�0�����y�ɓ5k�<��E�3t��IC�MM��yb ɑt�]����O�8�'	�;�y§�pGFtIԦ�(��d`���y�jE�I n�s �Q��` ��F��y2j��Д�Pk������L��yBĈ;�m+#�^��DmB�n���y©�mC ��.ү���Z� ��yRjˁ@���T��m�d�"��?�yR$8S-�a�$�׀'Ql�n8�y��>oU��֏����ub��Z�yA�o}
y�)_�n���B!�y2M�2���Ήj�ʨsש��D�݇��hP:�.)S5����pH%�ȓ6��L�n׻B�\�����VA�ȓs~�pO�<����'�>Z ���ȓBq�C�B�zM)�[9dS�|�ȓ��СR�_y�U���J�IO�u�ȓ)|�iAi�$�\�U�^
"�d�ȓ5�Ȕ�o��{1��ÇɄ�`I��?D�)H�'�X�Z7��>��@��*�
hK� х)���PI��_�M�ȓE����!�S�'��(8���ctޠ�ȓ�DT��`^�eB�#j����0���e�	�h1��J�������+��C�!��l�QA,gq��`I�1ApC�i�!�����?/�qU*D�$ɔIM�6�}X�@�u/��QE&D�,1qC��t�a��dM��) �"D����_3e5�����5�}zrA�>�"E�"�4��Ղ�
P����u�4qBPl	4���d�>h��fOs�!�D	�@�$HG�*<�:�S`����!�dáN�v��$�FM����#v!��"��u;���<��:�$M�c�qO��	ӓLHI��#�Q�(]�m�#nP,��MCsg� ��q��BI%�|#%,TX�<1��X%WfQ�!�G�pc�A;&�TyR�����H���8��.D�NJ⃊���p���i�2 vi�W͖7
�d)�����y�x �b�x�L*ғn'1Oƌ�e�F��3Ð�8�rq�T
O>7�'#]�9��!6`�j�jbME)F�'̜��D\6'`Nmp⥑�<�ʉ��Ş8���u�\)��($٤��4��{�&���iI�I|8�@����r��ǐ�<"���"���?��	��CQ��4aЯb\D"�G
/QzC�I�S�"�����pwd�B$Ŏ�8�"=��	�x�s  ]�C��@��n�M���ȓ	,.i��KR�J�|*fD%v���ȓ�t�s3��`�	�M���
E�ȓ��| q�Y 85��BB)Ҩi왇ȓw���q\ ?��A�E[%��q'��G{������`i���*�+:�p	���y���8c|���僐c,�yE���y�`Pk��!GFߧJ�������p?�O�چ	�u���
sGH!L�`Ł�"O����*�"_Op	��*WڢI���'���Ȣ*X(d�Y[g���rP���B!D��[f�Fuzd��f�VY�b(#� ���OJ���<���ǉK �|ɦ�	? �y:"�|h<Yb�R�X_�	�Ƅ�v�FA��h��ƣ]��Z�mO��`�B����C�az�R�\�'���9C(Q�[�g��-�8��	�'M���p���|fbm7R (��a[	�'U�QZrj���HQ8�ut�9	�'f�y�L�9&}�I���j���'�f-+�АE-�`�L��d�*��'&��Qs Ͷ�9A$+Ɵ*�<�j�}��'y6eb&���+�VlKBAQ�v@-��'����u�\#>��`�q�D'ox�e��'6��f��#��X��F�
T�)�'/dP:'�^FȩUM��~�0���'� (�i��M�*���D�=�����'��� )Q|��F��~�`_���B�ə$����1���#A�pr&��Y�B� }����.�2���K\�Q�8C�I]��  �Y�Pyj FЄE5�"<�ϓ0�8�!eG�F� �֏E�vj��[	��Ia�0Ow~@�f���1,8|�'��~҅*u���D̝<LP3&)���O~����?��q!l�K�$) �b�<A�,�9}\�;u���P�LM�Et�<�hF����oWP,�i����o�<��nG4�����3�0Z��m�<	���9v�.`�fg�*�d��ZI�1Oj�=�|R�bI-ck �eN�,v9��'g��:�S�'"�*�#c�-n�Z��@�_�E�����X��X�Rg��:)2pH�.H!M��%�ȓ]+ )(�m)�ΰ�S�SS�4F{���Ǧ�T��%>P8�	���N�`-���+D�$��V�$,���X�8Rb��I>!��0P����wb�)�������!/!�D�.	�^|��.J[�v��ӥ* L铟hO�B\:�n�:}v`uX���#��H��IP�O�p�b�ϕ�%~ޔ'��Z�z��';��C�'�	� �W)́s����'��mVo�v�FМy��`��'��\�sc
]��@��٦q���f�>��|����5sqVH�a�ۥ5��4���#(�!�Ow<I�@
R6�|AJ�LѤ��d,�O(�� ��&pA��p"�	7a�R	x�IN�OM�z"���~�YI	sLz�
�'y���&
P
y3��Ǎ�+Vܘ M>����� �A'P�k���+��B�X�q'"Oܹ9���kg�@�1�̝(�h��"�D=LOt���χ�z���E� ,7�L��5OtiH!+W)_���d�j)�k2��Th<�"fGi\(Õ�P� )��ӡ�OX���ܴ�'А�%��M�,�J��w���}��'��3ڙ?5��h�E 8�T��y"�/�Ş%^�]ʄl�F�Vh`�@�7������o������-$=�Ȇ�g���{3�	(x��[��3�"	��&�(ak���64���TH�d�C�ɩH��Y�m�3Y�Y �PB�C�IW#����
m��jF"y��y(�\����� s J8��!E�5�>��gV�:Z��	g����-��|�*�.�#v� ���6<O2�Ix��PU:!ͅBn��r���Z#2C�	�a%���"P?g����-<^C�ɘ��M`�\�bM���$�݌q�&C�I�kWp(��LS�y�K1m��D'6��E{J~�s�B�Yb���H�5y�6��F��!>u!��v�X�˥��U�dP!�"�; !���G�蹡$�4˴��a�!�M�6Ԅ1@��\�}��L�玖�}���>i������IR�%��*�+�"���@�E�!�$��
��B� �]��}q� ��$^��:�O�!���(]���
�h�$"O�UaR@�A��Ʈ�~
�MB1"O0��aVO�P!�5��[�h��F"OԜ�`��:t�I �A6i�K^��y2�	�%������"\f21�#D+�y�aԽW�Ƅ	��	�X��+�Z3�y�$G�2�\���o_�Jr�ZsaU �y��Y�bRA�u ��I!z}�#)܉�yb�Ȼw��� ���s.��y"o�d��=���$:������y�I[���
�K����SÁ��ynV6�e��'��3ć���?i����DŘ��E���-�w��w����FR��+ ╍H��K�NT�b�6	�'[a~rD�����O]GKj�S'� �O��=�O�4j7O urt�����"��(�'좼�c�B�.��\�eI�	�b$ˋ��8<O|�a��D%N؁�����d��""OB$�!�M	B!X A58��� �M"_Rl�=E���"hAC�� m��V
�"�0=�#Ȯ�l�'1�����%�t��ЉT���	�'r��b��{Y�;U��/K�T���{��)�	��o��%9��.:)��k��[�G�!��T�I��.*[���Ԇ�;��'�ўb?Y�q��;Xm�����'����'0D�T!�Z=}�Z@�c]�T�>©�<��'�a{b��"cGj����v�ty�$�ޒ��>I�O���H��d�alߋU�����@ ��x���)�#0�K0X����7��O����<�M|"�j׎;�b�2+�2I��Q��~�<A�D�
+�v�Ѓ攀.��1��$D�'N�y2d�	WTF8���H��Ir�Z�y��0&��r*U�GF��r�&�y��'�r(p�@�?��<��hћ�y�ĝ)'I��21��k3�aq��y"D�oI~��/�a]z���C���yÒ4l}�p1�G� P7@T� O��yBmOt->}s�A/L��D�g׺�y�]�G��g��~��Ǆ�y
� B�a�� Q�&����/�l�B""O�h��M�P���0j�XB"O�$��̀]��p�B�õ�n�qF"O��(��'�j��D�"��2&"Oā�*�2��ԑ�M�1P��R�"O�I�t��d�t�H��]8?���"O��$��|���i�3C�P!"O���W͂/�p��J\)
 #�"O��s�E��RdꁀzX�x��λ�yB�/+d&$9qD��lX�9(0��y���*k�h�ϒ����͐��y�%	�
$�`I�G�9��,���y��{��i�Vd�+?����ծ�y���6J�CǍ7�]ba�;�y��W\HKn���Q����r!0L��,�b�<�Y҅ުYH|�ȓPjyc$@�6�P��oZ���u��3R�e:a�^
`Q$�JQ-";��R6D4�C�8\F �4��Q3V4��I�z�"�
�� ՘LP�ˎv� ���HjD�0�T0��/�8i �8�ȓK(���ʟ�b&Ta!�MZ�nt�d��~5���ɦX���(ֈʭM��E�ȓZ�B���)�b݉f���B� ����"EH���0pV�q��H#xs�[��_�.B�I%,A(�k��L#��];�B���C�9I���31I��� ��G%C"c��C�	�@ÎXy��\�/�
|� �!W��C䉧<���;Pd��w�m��OEefC�I(i�����锅<ڸ\c0G�[izC�	�%�@%�B��89XIJu�M�3��B�I=6�I�픛s�����H��|B�ɂԺ@���2�,q�����c�RB�	�Re<;q�~!P|1eJh}
B��e
�|6�A� %�A���	�T$C䉡>�>IW�ڥd�,t�I"O %җ�D<' %�5��$P"O���f Ր3�c$�Q�i�LMj�"OdD�E�
5-D�b&b@!�Bukw"O�i�
L3ֶ@R��L�����"O0eÅ$��nc��h���9t��i"O�A�3�̺J8��E��5u{(0�"O*�J'`*]Av	D�
H{|�9�"ORD�K�H�r�ă��XkP�jT"O ���+�� E#c~:�u"O�\�T ���J�c��ȵ�d"O��	҄`�.�+�hD8.�� @�"O��ٗղ�n�`� a�\�1v"O aG(X���B�
J�&��"O���ϹQ	��"kD"!҂�1s"Oj���J��j�"�C�ڐ/�`z�"O*P{��*2�ꉻ��.��%�"O�`NYkO`�Pc�%z�js"O�p!oČ�b�C�'T�e�D"OT!���.P*PL+�+�����C"Ol�w��/@Hɣ���N��iAa"O��t49�aڣ���j��"O�q�\�5N>�:�HG�}����"O��x�%�� a��M�c��K�"O�Æ��K�Y�Ь.p8@�"OhG�GHZ5e
Ηa�x�"O�AjWF�6\����qIי.V̜�]���5DLM�S�O�<�q��B�J�T�k�iL�'O:�Z	�'�p �fԶb���e� ̀�iI��K�g�8az
� �� ��G�j0�br/�e���'�,�0Rc�	l��6���d�x�!�Ä.�L��ȓb�l8+6	�_3���C�>� �F}�+F1e��E�t텡{J^=��'�n��Wɍ�y�lԬ}�L��L�̍�U��~b�J�S��l�=E���#D�r\ 6��G��� @Q8�y���ļ(�ߙn��B�T����?1��r�'\l������yb0�f�Bv,�����T��q�L�(�r�2����5`�h�w�!�$[�2�(Ɉ�'	�b�҅����>h�!�ѕ8V�����I*t�)0����O�!�D�.!���G�X�s����V��OC!��Ky.P�%�I<v�(���Ŝ9_!�U�Q����!lF�R��ZG�8M/!�d�;��QRǔ"2T��Q���c!�,	i̩ ���j�����(TtF����<���,R@�R�WXH�f3Oh\yp5ɘ'���!6c����b$Z�8
�'���I�G�-s<��"���b�LbI��	 %÷qO��y8Ua��q�����KM�����"O((�Ҏ�;1��Q*��O�n�h�W�$��L���Ó���HO�1F< D!D.�\g�Їo�f41l�"^Ш�@�Ul� �u퀱� C�	2��xH7 љ;�j5I�����d��G`����y���tR�	C��"d\�$���yr�ϖ[\0�Bc�?(c媣�����~S�0ڍ�����114�9� $9P�ICeP��yB�E�Gƴ}:'�X9$�,=����=�yBl�w(D��.@!�B�KB���yB�R �Aw�Q"B�)��.ï�yRG��0���Lԍ�l���/v��0:��<9c���!a�U���}�(�ڱd�R�<�"I�Y�6D���]�[)��'��(��ݣe-c�>��QkE?����O��p�
e>u ��'l�ܨ{	�3�.�0 �3}��͸>�<h�`	�RH�R�Y�I�'�VX�mY���Ϙ'N�Jq#��0b���ƿ+����yBI=,���=�D�_�K�`y� � �8�*�4!�]��ԑnh�0rKS�0�arJΩ��٩�	�%]č�F�U���=���QwF�+T�ϯIR<	��i�V�H�w#��*�]$Py���q���'�~8��A^M�<a��S�F����޴�M��㓨LR���tC�02��ґ̖�{?1��<�X�����D�lD�aJ='�zM���'��y@�� ʆ'�+�qk�m�6%$����o}����	�5�F}2��=)Ǧ+��j��@���=�"m@� "�2`AJ��ydK�,�0����f�����D�@������d"����B%0�"�Q��OVp:�J�!q9b���Ƅ(6#J�ZH|
�o
�/m�E�s�� v��d@O�ɹ@<�0���'f�t�A,��!X�y$�,�7f�%6�
!H@�B�ݳg���(��$�7&&20*Y�ՠȄ7�H�������EeH<A��ϊY�H�3Ε,�����MKq��y�ԙb�Ł���)���T���
�i}B��ߥ� �Y�t��P�K0�R8&��L�����E�cER���ٓc������3VgH�!�m+x +f/^:�3��a�Rҧ��(���ؓz0��p�	
μ��D���DJ�)�q�O��|Y3��� j�U�s�U�Be��O�� gW<(�����zy �Ô�4�E�%�J+d� ���Q�!<@MY�>I��IY>3��Q D��zYTx1��`��Eۡb��j�t��'��9!~Ӳ�2O��	�Θ���"0��m�(���Ca�<!` ?o�bҧ���A�|F���ǅE7��̹����=a�M�m��Å�aӔȓ�����K��ûAnDL�E�ix���`Ѿg��dXX�"~nZ<�@������ �O��O�V� م)�)tF�
"��,ôa`5*�K�Ĺ@�k8d$�?�L�K�W�r ��񄂾`��9�v��&Ux�b�
b�"�[�*�0nРe�O6�|Ra�S��LepF��%C���ӌoj,\���׆�x�)W�o96(�؀lҲЃ�(I��?�֣��d��-�fm+?����@�v�֝�>�f�r3��G�6;����a�R��DS0l4�#6��?�b� ��Yg��B���k����Y���+���\?��ߋMgt�JO>��2��'����d
�!Ǡ����X�nZe���ë��[�IT�NF�I�M|"�
S�9ݨ�ZIʝ+D�=)�*\�!1�A�O��[ �^A`���
2���xĄ�8.��eDȹ0���0SJ\�FIԕ�ro-QG�ԟ5i7^>�cJ�1�69x5��:W�Q�"��hr��ӂV�!��'.������$� �eGQ��L�aj ��1�X�鄥<{�f�ـ�>}�'x��Xv��*r�<�+aIj�24���7��iТ���p�š  ��G1h-��b "!�ߜ����=C�S�Of�����c}�D"a�N1L��4���䏐/���Xv�%��'#Y\�X�<��""��Q��`y��>y��[�
���=O��U!W��h!�ɏ(؄I�D�O�<@�EFpP�N��YH|�i��2��q�ߥ8�ت UvDp�8�i��˓�0>���A�)�'K'8������_}bn��X64�9��|
���Ů	�%�س%�<��O��q�Wi��_"�u�kB�C�p�H�X�z��yζ���F��u������\�N�y����n�m[g*Z0y���Xy���� ~ļ�"�؃\Ƞ���(.�O�1j��<�
�1�
ʡaD�>]Z�킒	� ��V9^�ܜ[�<��42����f\"��"W�zH��KڞP�ܡ t�Кz��)b�ǅI���!���
C�
��g\b��MC�
�����TĆW�5�`'� !0��@ �8$�P�VbW51������enȣ`o_�n&~E;s�	\�XHFƽ��Q�'i�O��`�E#ɀE�������:"�'��@J ��|=QD.��3�X�0MUeJ��@�p�j5��jE0�V7��O*�=�|*�h�B"���Ս��h �%m�^̓i(�8Um��g��iaT�:]�(��Ʊ�@M�O��!�H7dA��R�"� ;4pS
�'d�ق�Ll�yPUa9zC�a��A�(�lm�T�S��G�Z7f��|��Z��y��#�B�Ո��H�0xib	ĕ�M��4�p?9B�����Y�0��I�3�����K\���t�?_�I�p-�ޟp��g^��=�O6��#��?y4��A%] A2% <O6�0�'X 1�A�t2:�`��5�XRF��:�,`	CG�PKN\	ش�M{#�$Y��J��f,��Hc�@+�J"[4$	�'�($�'Z24!�'�-(�(@�F��la���`{���Ct��4�.t��̎[�p �D�則3:l7툸 �8���' �X���U���!�1��4�S�O�}�F�a� TtT������
9*��il�v�;�n����L�B��rm �i�Դ�ߴ^�~b�_�Nw ��+G�Hp0�&@��Yi�1�G@�j$�!DFk.��V��E#Q�!3��0��,ʉW��q@���<�2"�Tx��A�	� ����B�(Ȭ� �3�P`Y"��&���;Ԡ���1��,�O����|}®�e)�3}�
��h���ض:Vi� T��'8Py�v�Tv�� �� kY�e�;��(��ɑ$���t��dD�3|�]�'d�����p=q��I�F8�f.��i��9�c̘�5�"��Tn�1n��h��
��9Ŏ�bÍ��?=�'W��!VLw����?v�[�՛M>�t��/4D�H# �^�ن���,,f�IW�Ҵ��ٰ��Y���"�֟tT(I+0 ^ߊ�m�Z?AW�O�M����}$΁���%;�f�G�'!��2i�&[F��v�BXԐrhS�z�A�!aZ���aM� �*��l>U�I��O��ʘ�Vhj�NM.Pni��$T�Z�F�Q��\�b�^A��4un~���
5�X�ݰ1�Ƭ���TS��e8UE�+Y���	D؟ �'��%x�C�f�f|��M or�@�G��0�$�\�0��������yw
�5|�!j ��3p�L��ƴ�y�A�50Y��Np������{Jucc��r�t7[���OBĹ�}BK���`* �P�bt`�� 6�y�!�=NPu��[�AдԲ��̑�?ɳ�ՅXv�M"T+lOԅ#qj�"(��M3N�����I�u��ah�Qz�%#��7-�7c�	�"J1�rU�B�^qJ!���w�p4�UgG�Ȗ �����E'1O���퀮F �MJ�Is�O!���dH*��|P���61���K	�'�)�`Y �����B�)a��٪C!�r�U"����E�<�F"�i�p�[p�Q�u6^�Y�T^�<�4i�"� ���B��Q<��C��\?&a�'(�����G% ��k�6범aR���a|��LS��5T̴[�@ '�`��F��|!�ď +Y�Ej7��/���O�Yd!��R����*��BB��+@b�!���?�
�PQB		3�ٸ�-ߙ;�Q�����'�<�[�+N�ܱ���T,e�����'@*�APN�^!#���m�8�bݴ?	�-�Ӏ��dea|
� �a2�/Y�s5��ue̚
��0"OT9�1��Xq��)w�"0��"O. 
Q癣8ɠyy2!>�x�a�"O���� ��J
9aՖ}?�-�!"O>E�E�'.l�a�	-8���7"OP��$Z��r��f�zDCt"Oܔ�V�Lz:6КSOA�q����"O��[��
8���1`-V�<(�"Obe8@f/��Yၯ߈HԬ�a"O�Ih��_Ղq�"$T/_j�T�"O��Jf��fg|$DÛ-[DEG"O^��!��	@Z�P��6O��xc"O�,��k�+�����B3����1"O�P3&LP��L���[�4inE�`"OTT�u��<#���_�7����"OJ����gN�	�pl֓ksB�"O�L���;X�|e�r�
j����"O�����Q<U�%I�
��!�D	+�"O|�`��NW	�QS�k	�T�8@h"Oʙ�`��(t����I�
���R"O6��WE�0������x�@)8�"Ov �B�Xq!��e��W�R�"OU+�A�M�:p�w`ݔVE	"O�X�"�߭.-zqR�Oӯe(ltJ�"O�ȹ��߿1��e��}�́�"OX`a$l��m�B}Hv��A��P��"O���P]0�a�&��.�zc"O��:Bk�$%�4eȔ�S����`"O��XA��v<��!��:8�ڠIw"O��j�/�!`d)����H�"O�0��J���*�X�&ͅfҪ� "O��Ka԰�0HXP�^ t���T"O���@��)%���X$�ˇ4���`"O���kS�݆��%K7T̢!"O��)Ss��fI>9h��i1���a�!�$��n�����F�Mr��Dw�!���'~)�e�1ǗB�B�bT�7&"!�D�^et�Ɇ��Y�PT̓-x!��ޜ"�T��u�ߕ>q�l�6
̬?7!�d�O8BQ2MY:д@WIK�w!�Ě�*��q
#��%~�,U��i͑-�!��̖w����q���g=\I��h��!��2[��Fh�w"Bx �B�{�!򤍴N�����k"xc�Mé;�!�P��x#��ɷQ,`��=E�!��|��I�E ��s�Ċ�!��4oZ���[����c�\!�!�䙨S�^�UY�p�*ƀ�&;�!�j�
�ش��,�t��1�S�,�!��ѼNJ,�G.CY���q3�Z4�!��_8&%t�Dᐮi>�H4`Y5:�!��M��Q���5q�&8zA�Ҫ>S!�D.�\����\pț���jG!�$C�]h�����)&�hkơ��&!�')M�d2�b@�������#C�!��E�ux��ƯY6Z�)�F�]�t�!�OO^]���*4���T��0�!��C32B�!j5mŊ���̏m�!�ң$Ϟ`���m� �y��^0Ar!�D۬o���3S쌷��d"��=wh!�dNZ��!rBX�ny����K:w!�ě6T�!�pn]�d�T	����e�!�dҡC���9ūC[�<��
�_�!�dԿz(2���ZH�Y2��2?_!�� ���wO�0����ß�B�*�"O�5��+���� �#-�|���"O`<A�.η>t���Q�r+�$y�"O�p���ϙZ�4[�NAw~5�"O�P�*�21��� �l�{l���A"OA�`NT�6!�@�C�(nV}(�"O�q�K�<��<1W���F"O�I#��70b���$̦_�|���"OtA ����9��� &��
c�5��"OE@c&AhlT���62��*�"O޵X �G��!�w@�44�s"O*�q��.[v��P�n5.q7"O>B�
/E&�´hÊY':1��"OD`�w�.`�d�r&S�$��"O
j��	��T��+P��f�QC"O��S���#nf�����QpX��e"O��A	8)V�2���XB��"O �]�<�,�
�
.< ��D"O�H�e
��/0���ʚ5!�0Y��"O�����[�}�Dy�"��G����"O���hO$1��9�MT {���"Oњ��J�`���(f~p�$"O��!!�49�*��`�С+D�Q�"O�)0�ּ��� !L�"�2�d"O����(�h�qRKF"��u"O
T²��.p��l�=��"O���KK�^�&��Ǣ�o�t�"O -�d˖1DA�=�D'�ZG�u`�"O�����Z����;1�+P�R�"O�`q�?��9 $-�3OY5��"O�9;�')6�|@��,Dj�ع "O�`Y'�7�� ��[�
0m�A"O�I �F�6*N"$�ƃ�>n�Y�"O*l��6F v��Ej�.p6�B7"O� �3�T�"���3�կIxl5��"O��QHR�"֥��D�mnB�Â"O�f�U�}��b��� 1^pYI�>��Dݑ `���?���&4�={�P��:D��)�Q2|@6�WLD58�Δ��E^�	59�Ā��8�3�I�b�����R5�f��G茟%�.��$��2|����hU��
��	H�((���+Zf�lj!��,BȜ���� (�`'gٮ ��f�_�x���POC�c;@`AO�X7pI|*� Sg��	�K��_8Lq6nH�<!í��_�@e�D��&*���EF�53�V����7I3\�bj
!^f�]G��'��<�fcB�pʀ�b�w����
�'�(�O7��-��i]9a��P�	��,��!���ؽsa��F}a\�M4X�Z���A�<)�e���=	$/�\*ԑ#W�ܮKN.�+�	}�<�C�7B�f�&d�?����DJ=7 �]��`܎Qq���Q#��O64RBW�|dN����@���4�K|��װ"��Eg\�!/�P:#&Gg≸9AZ$�d�'��9C���+�vjÏ#�|��3�14����W 5�&(����(�~��3��2������4Q��0�`��CA.$�\����ȩ�m��s�r�fd�զ�C�<_��0Q/Cӄ���7:���E:}�;>��4b0��z6	Z���QIl�C�%ޤE(�$��6��<r �ܱ�,,�b��>ƶ�J���#�� HB.�.�C�[j��ә~�v�����`4L��G�^�p"<���U1���x��	�v��h1ckF��aKǍR:*9�IB$�y�V��$vV�x��h�ࡓ���v^TJiS7M:HC�F��8K��'>M�mÐ�
��E�J'���"
��I��\���C(]�𤗬"��1ZTmCs00| T�% 2��A�"�qg�CG}�떐t�=�fA{�4�L�R�&�y�z<�&�
�D��;G�' ���a�v�F�n..�RTQ���y��,���|�t��'.�h���L�L��S�O�&%kv�#H����
OK������p~�}�LNs�O!�°�Ս��y�"�	B��`��O��� �ʨ�����S�? ԝ�!�ؾ>뜬P�����nl�S�8��ݻ�nIJ��4�'M~F�W��S*��1� y�FQ#H:X�y	�'��d:1\?%5�䱄I�?�V-A��G���NH�@�L'���'�'�iݹy�@ƕb_�\�
B;X:! Ё#|O"��ţу2�i� F�9b �����	`16�j�̈!�$l��'_J���{�S�O�0�h3�Z�_�kAAG�2�@�ш�d�(=$u(��4Z�8)����-*�@�g��y6~EAB��ēY�d�҆��p<�U隙0�����κ\��5IR�R$\���C��`C5�ݯDŘ�)�'
�(��-L�\z�����Ui�y��˒6/�4����'�L3 -� ]E��0 ߨb�n)�q�.}B���U����cD�i�Z �	4��O�d��*)���ڱ˛.6"�����p?���!���cuA�3YV��x���Ya}�3�C�U�=�5���Qs�`�E�1}���F��	f+��L2�jUeB9V�Q�Lh`�g�����	4�����+zly5��
	��_Rܸꉋ����. �`�A��9Y�5��)7���ȎY=��
@M	���)擩5�4�b�Z�1���A�D�4�*D�-ز(y�	B1OU(1�H'xbx�L�==�,�iV�>�rŘ�~p�y:��ʣ!J9��M-S�ӧ
e�H���['�Hu�t۩y]"��D�
�Ѧ��r�<����1R��5��@�|�ٳ!GK#9���l���)�'��	�� R�pRp%�p�=D~R��b�
�����J�|�tm��iyȍ㫋��'���3qfWx,�x��O��4�G�1��ÁE����DP���hh�/'��/W�:!�W�O� -cv(�9px���"��x��N"ZtRy�����y�Z�	�i8\��'�^�!��9ݘϘ'�0H3�ұ7(���Rc�0f���
�� �(p�޵6
�b j^���[DI�$��ECs� �O�#��]g� E	ED��6�����/uo�)Ӵ%�h�O�8���T���aR΁!U�6��	�'Ƙ� ��W[X���(E1@�h)Oh!X��Ӡ3�4M��|�1�U�Y�ȹ����:i7!bqg H�<qc�G�z���[5�L� �ҿ5d�k=�!���'��g�h�W[0p�Ȝ3�l� v��H�'ê�Z��(>����N��0��r��$t�V�ےßi؟4i�A��U���*X���
��%��$WE���5�d�h���[6AǸ�jg��)"�2��"O�)#G�ęm������IsY�P$/ϑ4txӧ�>E�t�E%UX�1�"����ѐ�y�Y�	l [@��5�����?��'��Q!����Ϙ'��\J4�	A��`��a	�!�'A*-����:�jH$���U�X�ȆΕ�:x�F4Rtp2,�	�0"b�T�Q��E��
�|(k��Z�H��@����R]��r,*�/]�$�pgŮ�Gy2L1 p(F�D.8I��Ux�Ɇ�ݑ�Ǖ8�y��_�P,�'=:*�v@|��E2Qe�zɧ����er�n�U��E+]E2!���q�"\r&]<;�2�9Dl�%j��k�"`�ك�k�_؞�82雱
��X(�CԢj�P�(16|O@=�K��Kl�(ڴ`���#��L�|+d�?W�݆ȓi)��� _�j���z�g@5%i���?���M<V�J��!ҧ�n�I��XB�͐J5��>D�P��[1Y�đc'�6��Q� G�=��)�\8��N��~B*�/Qz$�`vE�Z��8XI��y"(�j�*m"(�X�R�Q����?�FJR$T�`�j%lO�l0�B�A�(ݫ���x�T0�'O�����'ՠdlZ%T�y��.�-Ʉ 0���BB䉊!(����A�YW� x3�-n���أ���D\�#�m{�𗏘����`Ã�E"O~]㥡�"ck�GV�f8t��W5\@<�&;��s�@S��_� d0� 5�5L��tA8D��/4ؠp'��7O7"�ra����&�8h]a|ҁ�(���hu��(��e�C��y�[!�Xeb��	]<Z��.�y���|x*��"�!?:HK�C���y
� B-AV�3>E���'� �U"O��H��G��&]��ԗ~��=�"O����iV6��X 4#�f�2��F"O$�I!�V�z'���,�x4P"O��rԡ�6X:�sb���@���"OQ�'��t�H�A��ɚ�"O�i��|xNHY'/C�Q�*m�"OBD�e�ѷJ�NH(ql�GW �'"O���H�>?(j��)=\����'L�)��@\��� "�ޜ��'�����n�n6��;�f� �����'Ěy�6�� �
�:��T8�>�+�'��7@�#$�0�䥍�ozT��'�P�	G!Í8�\�I��xϐ��'���T(7,���z�@5{6B� �'<ls��4jh����Ǽ}�\�@�'f�h��ʖ7Y^81��$��\U0�j�'>"eY$iL�{��L��Q���'�Q��l��[�����c��S����' +�N�D��t��G>C�	�n�E�U��-� �����6B�I0v��1��aNGj�Q�B��A�C�I<FR���Y�D��vΙ��PB�	��b�3(+tR�|����2
B䉯&�9yW��?hj<1qK	n8ZC�d$�ei���5"9�d�&*��B�	=4��H�=h���EV`�B�I�L!��Rq�#Y��0&�VI�lC�I0�2���Wj��tc˺u|C��(f�&4q��E����Ņ/a"^C�I��]���><���d3/!vC�3x3�dc@�iı
b��P2��$̫����QG_~}����,X�8�B���<�!�v���oOJ�$�!�?�!��5�`e�l��Zj�������!�Y�`�*����LH�y��A8z�!�$�9J��A�ʱ��%�2̌��!��<�|0��锠>��\x���6�!�4\WJX:Ц��T�ڀi�*^�!��$y��8x� �	����cF�4Z	!������q�Շ_�	SP��95Q!���#��<ʱj�	Od9�6�K�!�D��~k�t`�͆I$hJ���o!�DӸg���O�&�jt�GG3dc!�&����Q�5,�#�E�o^qO�FxB�b�q�(O�$���vF�	�BW(��%T��a�3
rX�L<E�d���\p'D&*����NQ�?����w�B`�B-������,S��Ku̘5V2�w�F���:�ʀ<TƎ7& ����|:��,�Qӈ�?-A#�����蜤C݄��d���4�Rl��`��M2�mȌNg�#n�	U���k�Hu�d��(Ăq��X%�[8&�%Y'k� ;�@( 9��غ�*�
~:&Y�P��(A�9����-;�@��Cҥtn����#�a����X��P��X�Dw��!DB9*��䁥��5ʊ�@d�ښC&��
ç`���k��Y���:I%6P&j	:�M�0�<<6�I7�������s�xXbk� �K\
�XmRci�+&�(�%'���
�ZiZsI�O?��?��MkV:"�.%�f�ӗL@��sN�4fd��+b�hw�)�x�O��+b,_�NѾ\h��ֵ� Ԙ�N�9"��c�А��?���(����a"�Gkc�a[�)���'�4!��S46}HcR��"����ݱs9LC�I����a����>��d�F�;�C��'05t�d�ƉD��̈W���<�C�Ii ��B�G�ޜ���P��C�I�!���4�t�N2$|.C�ɏ.�X�+p`K0�60Kv�9�C䉢_��;��"F(t[5��/@ߌC�)� �и��(4��򥠔:%�U[�"O��%
R�AS2�J��3cf
X�"O��[v�� 
�t1q�!�"X���"Ov\1�D��u�tD����}���� "O6��U�%h�`��O�{X��E"O&dѡ#�*ޖ�{GW�%vtH�#"O
)zT�KY�ɳa��$�ha"O�\�D�:N%����M���l��t"OX�2����9�\$�FlڠC��"O��NK�6xj���J�5E䱊�"OΘ;���X��K�GטBJ\u"O,��q�N�F�rt���R!2L,�R&"O�$�c��
\)Dɘ4����"OИ:�@�4*r-���Z�2Ep"O a j�=IF4�b.�2���'"O摂��O�R�}@���5N����G"O���K��UU �(Aa�L��U"O�Ա��e�	�/��k��$�!"OrQ���~d���t��6�J�Kw"O܁�F��)oV@LR�+�.m} �3�"O~|q�'B,M���P�+�-x<�t"O���ǥ��:��p�_�tg�eش"O�h��T��<\����	d-+�"O��b�E�v��c"�ʌv�\�"O��$��E���qØ4H�l�ۆ"O�h��m�7پ�����8�a�"O�4���~�~Y#b�^�E��"O��@D��!o�\`#��"}�es�"OT�Çi��/h��� �C5����"O�-(V'M.~q���1%֌��"O��	Kħ�!qt�*�S�"O���&�Cg�f4P�CF�Zt� "OȔR�� �4���A _[[�u�"Op��I�q�H ��Ό_Y�X�2"O��V=q>���M�:= �(B"O�i�S�!l�.�����([�F�cE"O�a�I��b��˩s�kU"O�4:�����8S.ƛYx�2"O�9�a��^�R	"ԧ�8E9*�"O�蒂 %!�� Z �-<�$�%"Ob����F�iV��"�-0���"O�P&��	$�1"R;I"��Bd"O�@��ǃ�!Y&]KB"�
PtY "OvA�i��u�l{��<+�e��'�8�kF)fY̑0.Y9'�RLa�'�Z���-F$JP(!"]~�#�'o�����Ə	��q�I�%���'�Ƀ� \;	.B��3fV�f�
�'����n��\�FJ���GY��y��Y4f� �����P����y�.J�?��� Յ���BKH�y��#bz�5H��k �Q����y")�%"5Iq%�ày�/G��y�	�K����Ǒ$s5R�0�yR�ϐ,�sT&\s�<���5�y�?����`A�� �8�ؖm�3�y�LǕ�t�ܜD�&q����"=!�޲j��u*�^��RE�t��!�ě�c��a�j��o������5p!�D����{�@;b�~ȀVJ�F#!�d�/l0�u& 6��00�i�*
%!�$ӑ��� �ʽU�^�聨�:!�D�A�-bB���~Mc��X u%!�>yr��e�L�(�a��λk'!�� �ب6+̀� ��r�	��"O�)۷D�t��	S=h�V峥"Or48�G�1LpZ$�`��gݲ��d"O�U��쓈�,�q5`����P"O��ǌ��x��-�'F��X��"O�x�g�r���]?EPI""O4�f��$���!�ˠw�����"O"�"�Ŏ�(2����(>Z����#"O�xyŌC"
bL|;hM,3�l���"OGe��Wnh|�q,��%�`@*T"O��f��mN�{���
�F�� "O�)��-L�F�hh)��tv.�Q�"O�%-)Ad�#��U�ge���"O��Am�j|I����9h@~��"Oz��b�&P6�u��%E6r(Z�"O�x��,�*4K�}`�억uv��	f"O���P�T�� ���[6Rb�� �"O���Ń��j�8��@	�=nO�)�v"O�)�ϝ&` ��a�m�I� ��v"Oؤ��͂j�<`8t�k64#C"O\ucQ�Su*m�E@�d�9Zc"Oʑ���>�pA�Q�г�"OV-k#,9�v!�)�� j�1�'"O�u��JT�_�1�4(c j"O�q���{��!��E����P�"O�}��̉6�h�Yօ�?����B"O�Eyr�	S@nTx�䙥l� m*�"Oмyc�>d�Tt;�D�>uLHI'"Oyc������p�!u"O~���"fV���ڪn��("O����$I�E
��������T��"O��RH�'���r�aÃM���b�"OT�㘽&�\8@�NBud����"OlE���[;f��i� O�~��̢�"O�t����(�x�CW ���!�"O`���Z�mh�LQ��߼�4e��"O$���j�$@����4%̙l��QV"O\�
|������0-�"OJ��d����)iC�4?��Jw"O�\��
�%	�qe!�2�y3E"O��еMM27"6�X�)��P�n�""O�9�q�M8K��(���5� @[�"O�� �L�5hn0����6{�p�"O|i�p�[�m~�i����rL!�V"O������n�p'�S%h�@]�"Ozpjc�"S�;BU:� eX�"OA�P�*Y��N�2�AP�"O�̹�w�,�Q�JJ�f�@�"O6􈆠�8��hQ�#�2��"O���A��b1 y� *K�D����"O����%D�
o�Q�Q�Qw���"O�1���o&����Q�РU"O@xs���R��rY����"Ol!t��mт��*��QLʝI�"OR�rjz���5PV��"O�R�֑D|�1�GP�A�"O
�Q�T:,�)Ȳ�Qm�6��t"O,a�F�̓X�L)��cC�5{���"OX�6aӧ{�:�;��$�"OJ	$*F>P����J�Ub�}��"O,��Wf`0Ua�Gny�@F"Ob�ơ�gzB��9~|$�G"O��S��8�L����MZ.�
�"O�D�$��	��0��K":Sb�H`"O� j��1M؁Sƴ% � �So�1y�"OB��AhD7(�S�)F+�p���"O�� %kD�9Y�4v(ȷr�䬉�"O���@�֤o\ʱG��Y4ndQ�"O�2�͚;:<`�R`·N�92"Ox:o�I���ťݥ<�&�R�"Oe�DV�ub�@ 䈣\��"Od͐!�C,V�.�2�b�4�d@�"O�]ѰN)LrH�Gޠn]"q��"O�A1��9&N��sF�2��1;�"O��S�ݤ"^�� %�D�Pe$D���q��{�xU`��iئ`K7#D�$ç,*C6���F0�4]pp�!D��2��N=N�a��5�P1��,D���'B�>���:�΃�HH^�Y�
-D�$jKF �D��+��%=�
�)D�H�jW� ��I��߫k���:�N)D�ԉ�CM!C�L
ǃ§*��U9Qe%D�|Q�陓
J�^�-$��KAk5D���A�a�<�C��^�����2D�(  a�b.�«A�8�p��"1D�٤폻Q�0 R%��z��$��-D� ��FX�^%��[�z؇���y�爬 v�8д�A�5�8ܰw �y2�<X'���0OD#>M\��.���yb*�6����!� 2��L# 
��y�̻%V�`��� <��Ʉ��y���>�I�cĂ2�4��"�$�y�V�-��DB�xo��2�W�y�9l���00��t�r!�jê�y�
):,[p	 $�lK����yR�	k�<���i��I�i 
��y���!_�d2r��07׬*@*	��y��"�t��.;'̒��yR��=>���I�&δ�&�;�yRJU���xŭ��f�n�jJ!�$H�)ڠ���'lO c���-!�$����y�g��N6�Cwƅ�n�!�O~�LD��K+0G��!�z�!�٨h��=��gQ>�>�jW7�!��8V~PHP�8:���� �L�}!�dXD\B���P	e�I+}!�ӑH�X=ٴKU�2�x�A`=v�!��קR(<��*N9���5"�>�!�d�ܘ���.x�� "äF�!�d 6��H�b���a��ķ!�!�DǍ��-��#� 3:>�Z��Әy�!��)�R�`CaQ�q�"�3a�Սh?!�dT��[@`D�dd F���!�V3/��b W:
l���GD�,i�!�$����B��&Eܬðcē<!�\{��"�N�O9�rc�&
�!�\2H~�����V!T,��`�!���~�������,�ڃaӴq�!��M�a��:��J���J+!���y^Ġ�׻s��̒pM�/!��W�/f�,��؍L>����'1`!򤅔2�pYT�ؤI=pTcp���ri!�Ǵz�ؐ����-�@��8R�!�D�++�``@N�6��X�"
	A�!�F8i�-K�J�L��m0HA�H�!�لg$ �  ��   �  V  �  �   �.  V<  J  �W  �e  vs  2�  ��  ��  ��  "�  ��  |�  ��  �  [�  ��  ��  q�  
�  z�  ��  Y�  � 5
 � � " n# ]* �0 C7 �A L �R k\ �d �k 8r zx �~ _  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf"O�Ya��=!l���Ɔ�b�V��!"O�!)��Y�fx���eE\z0	J�"O>��pg�0Z�2=�C�A�Hy�"Ob\B��;h�`��Ɇ*���S"O�h�T�ÕZ(jܫ� ��+�Ƚa""O�A���I�{"��qReM.v�\�J"O�I��cR�G�Fm+De����(�"Ov�M�{�Ҵ�U���F�T��"O� ��M�g��l�a��8{�Y*7"O�Z��іh��8`�tm�`�"O&ESS��M�,ɠ��b��b$"O,y0GD�!�<�Y#dYF��c"OV�Wc�6�:�3�	�C��:�"O�`y!�������3-�<�"O��!S��3C����ǇZ��\�C�'��	�;��0�Ѐ;xܰ�c�� �B�	�mi�i�OχF���)  K
!�B�	��:p ɥ%�HU�WJ<3��$'�����Ot�53Fm�(0�"X�vJ1D�� E�,]ʁy5��V/�� pK.D���O��B�H�#f�Q�f-��H�#9?��$,�03nE&��5��jF�H��	��'�% �H�p`|$� >�=�s`4�S��?� ac�Y���T�F ܆F	�g�l>�S�捈]9�0���_���+�������]đ�&��q	2��>V b7m=�S��M�ǧ'0����
I�(#�L�L�<�T�јL�4ě�1�*�"W�L}��'�UA0��)x��� O��S�l��'Ƅ�QQbY�O�z|7��H1&�:�'���ص�6O���6��M�x<�
��(OH�(v� �m�V�8Si?���9�"O��@J٦��Ui�hA8B��=����~���	B<(���0��D�|�,i ��
�'�l)���Xh�lY�SJ���
�'�(�4��y�� �˗�J�2�`
�'��A��Cb�>�)�ڈBS`,��'w���Щ�=P3���e�2	Y�`�'0Ё��q��ÌY�# � �@-D��@�@^�{�e����|��� �H'D��#0cʭfa8Kg'������h&D�̓@���[7�t�A�exE��,(D�h�"�,3�.Á:C��%D�B���4�"�2��4G@d�B
&D����Ϩ ��ؙr�د�`�r	0D����
��r��A�I�81 =�c-D��hݧEx�1!*Ƅ\�Q1S.*D�8�E��tn܈����;6�+���yBo�){��%KV�T�u��B��y⁙	B޶�TaԑH��`0n��y2�ݷ;v�}#�,ַ9���b�ǵ�yR�P�L��R b�3�����<�y�/���bt�Ra� $�����a �y���0]j\a���q�H��Ǝ���%�S�O� 8�ìF�UX���B
݇��D��W"�"A0�IF���\�ȓu��*sKH�u�h	+s�X�g��y�ȓuʒ���w�m���]�p���ȓi�Q�!�/e�@쑑M�'9e�P��w�ƍ��k�k�f5/�T�"d��J�<a�c@���i�⓱�.��2��I�<p%�@>����H�4�*��d~�<�1�ˤ#�"��ai�$u��@�
]w�<)DHK�?.Ԥ1���&'~
�(�co�<a�n��<�B��!�fa��(�h�<��(��;�%  �,���G\�<q�(ZRВhs$���}=
�S���T�<I�� W0�e��4�����N�<���).��	�K�-~6,�dc�J�<��ŌTD���W<6^Ԃ���k�<�Ѡ�;� h됭[Y`-1�`�<q�is�0u�|��!	V�<��
<�*�͂�dH�� �TO�<!�����:�-�@��9BJ�'�f�3a��'��1�Į?O*���'�vLv#��3r��QFĶ0:����'��h��l��CD�_�&�p�'b���+�K�]
wHȌ�@�
�'�ęO-Ei�xPv��w����'yT� $��}.�11
�4.qr���'��D�b�ϲmB�@�@ �X�P�'��D�S��<Zg��� L&� �'�D����"W��1���MF8Qh�'�h�gbZ%-m���K���a��'�yA���U<L!#��|ϐY�'���S�E6H���)�p�!�'B��H���!GBt��2(٢&��!��� �1�P��+��4¤���P95"O44�d�d쩠Cݦ�p�Q�"O��:"Dϊg�҄����{p��Q"O�eZ�B_�*;Ҭ #l��SI�Y��"O����d�� ��E��,��R#�'�R�'���'��'���'&��'��0J�%	!�n ���#�b=Hg�'@2�'���'1R�'���'���'�VD2B[�:�z��#@ʠ
�2U�5�'���'��'���'t��',��'�Z�ؓ�L�'����C�!�x���'2�'���'�2�'�r�'��'*Q�^�2����S��t���R2�'�b�'���'I�'�2�'�B�'��=;%��P�.\rCI�z�~�Y�'���'+b�'���'�b�'���'�T��F A�[���ӗ��+1��bf�';�'2R�'���'���'���'5<�0a��3X&�ڲ�	4x~ �f�'	B�'P��'���'��'r��'�a��.@."P�����Fp�u��'��'�R�'7b�'�b�'z��',So�T���Q���p��1Ӱ�'�"�'���'�B�'i��'r�'<d!��IM� ���FҀa���3�' 2�'Q2�'R�'(��'���'.
Ys��َrS6�A$�@o(K��'���'i��'�r�'EB�'eb�'�&8&FCiĖ|ـ�C��6�'��'r�'���'zr��'-"�'߬�[$�Y�"1�I�2dG�5�Eݮ�D�,��I��D�<�*O��OԀ���F="سeg@�V?�)%ˉ�;�z�X5���qڴ�?�G O��<���Oʭ�c��, �viϊ5J (Z�4�������k#~�\�2�����º���_�j��I.,�`�P&a�<V�h�ӎ���`��i��#CD�oe���'=�S/:g�S!h�v<��I3L7`�!Ez7X�$ƍ�A�b��+sU~����wLJ��W�'z� ���C�$s�=���'�P�j9P���M���9Ο"45�f�5a��%oT �%i߀2<�YSI"=�2E�^y��+3��O��ۓhKVy20O��+RB7���?Bfl�;#	+2U�m�%K
����<�N>Y�
C���<�b$�(4�X�6a�yR#��?)q
]|~�E�>)��?9q �.��߄N%d�rCbV *�`lIe�;Y�
�h���<�B�i���Zt�!���/�H9��'��}���D� �kј_�JE�B��=*�z��'b� �H��!���'��	7]�"!�ph��w�	�w�JZk��I� �~ �TF.?Q'�i4�+���O�P�t&��E! !1f��f�i��aQ�n�z�'v���T��*i8�NM0?����M�`mkݱ�fnO{�	ւK1�P��ʐv�}� S�Tp��L�"��6㕈�?!��?a��}H�,aC@Lw2����=_vpȒbKѲ���+N����&�O����O2�	L-�ʓ^J� (��y�8�sPh̑ M�Z$T��
�4'�������~�6�t<�O�&|y1&	SZШa�[�$��A8��N3JM�hB/�- @�iIs��`�D�����>1a.�O����W-/E�% ��D�)�x[dL	O�<�:��O:���O����O�˓P��Ő��D�?��m�3[��s�C� �J�"#���?Y��iz�"]�����@}�N}�H�mڬn��}#w�2� �H / ��OzXИ%�B�F���QB ib�;��f���0���B���M,__�h�N��;�%@Q�ZDV,��4N�B�'��O�L�1���w�0U��'���T��L���	f_�(��3G�&�fk>5���MK��'�y�e��M�4�
�!���剂~�����J?	�T�p�{��|2�b��u�R�}=��Y.�&��F�_�%q���ՆT��֥�A��?	��H0R������$�9L�ԐR��O��D�O�d?��� �����#G_$T����Oj�c��pEW��?���?��'iE����J%Ȟ���AX= �q��i~�N�>qA�i{v6MȲS]�dX�x3�O{�H�WlA.Z�)7�`�F�t~�%�7���_:�)p�L��y򧋤���I�
��1K��yǦ��j�z��W��L,1`[���6�'/��+�l$8����D�'�"P�@���e�,Q9��.O��(s�ʰg�N\�G��Uyr�xӌ�D�.5^�I0��D��I�&'�T�N̈1J��1jg@���Mæ���+���3���&`Γn>,�Q!�t�9����.��?-(��0�d�t�[�C=	��o��T�A�.]�6��	ڟ��I�?m�E�	I���5"h�B�E�^�4��X�� �U���8-Ot�d����6������]�G������"x8p#���X�tZ�4C~����,�~�&P)E H�OoVXB�����ݳ[J�����G���
֬�x��c��'�4��d����U���"��,ut��	�w��񰁖
Y�)���rgXa��֟����0�'g��*n�
���ԟ��Dg]�����=g-�<I��͟��J/?�^���484�Ư	�~�&�<Z_,����׹Tf���eC�nv�7��9�y�jS�l>Ux��=(�(���'���!6��ğ�{"�D��S nP�~�z̋Dń1x&�z��'�r�'�v̢�%ŀ!��O���'�R)]X�|`�H]#_ *AJ���&��SM�(���'2*n���[�u��i�]	�H��0HP�"�+Hlijs��<1񶠛��M35i��W)���[w�ʼRs5OF��%k��uF&=4��2 � (^0�%@I�Z�<`�S)��<��.�?a��9=)��9���?����BC�3lS�����/^��:����mb& /O yY�BٖT���$�O������y�9�����*ܴ�0�(G.xD���D��4��'yt7M��=�2ƣ�<UC	%P����+�@�H���|Qbt����6 Ҕ� ۀD��y�R$|������<���p`&�I�L����	��z5�с� !��jƊް0���{7J�'r`����@�	�4�	Ey�NF�#���8OJԋ%�Ĩ��g�J�y�" a�'^6M�O �1����8)O���c�$�0�f�9o��JtJ�h�9��#�p�J	��� {R��%��3O:N��$�K;f�H���+��S�hG� 
��gIŬ&��0�/�p|$��mP�	�V�I�K�Or�D�O�����|����R�����䬎�Y�Je#�K�*���O������%�t�<��i�r����y�[8�=Z�Sl���*Ӹ́#��eq�'Ĕ��5��^k��OW�!� ��P��o[�4���х�����12��4��	ȁ�'�1B��'wx�`$e��sr��P#�ꐋ�<Y�	�p���� P�f㍷L�xi���; ߖ��	�H�'�&�3R����'V��O.T��3��.�^���E0�}i��ݎ��I}�}��lZ�W���	�6"]q�;�=Ɖ̹ØQ�C o0�uc�(>�������6S�6O96�	��?�C5y&�4��@�S%қ`M(-���O��s�"�OZ!�d)P��B�d�O��O(�d�<A2��m-Ⴀ�c�\����:dbY��Y��������	�K�P�|��I�b��P8Kt01��kX�7�� �E�5�MSei�$
�X��I�=zX�+��qzNM��v�a2�]�H�ݤT+��3R�|��T�QF���IJE��O`@ІH�4�����O��������|��h�T�$��Uؾ�+f"�_0[����?a���?9��T�L�,O�lz������8^��SG[�*���#딼�?�۴}�H��|񾘊p�;"�C���uw�:�	A�VBf�����FE&i�8Oȁ�+�(�?��N�Q�d�BZ���Z�&���O�����ߕI��qIڿ>��4�U/�O����O��D�<�F�E?KWB�2���?i��#��T�@��=<2��2�zw|H#��ijĽ�'���Io���fӴA�O"�X��M�8N5;��8���g��Kq��:�'��,���
�OS0����1�yB(ӝG������3-Y �l�{ ���kY�)<p�J�=��'����A�� 9�����'���'��`�ڡ�*`�@ʈ>���`��'��"�EM��I%�M��R�A�y�h�:#yB��g�_-,urfCDg����c�+��7m��gj��w�ْ��P�<y���#��� ���"�i͐H�d����;mx�����
���9A����7���1��O����O��iX�^M�hb$�ʩ`���j^�Q���<yv��O� �P���?����*��_9���32���;��͸����U�G�z��'/�7�˦�蕩��İ#����,J̈́Y@c�]�:��2uFF,��IN8 Ly$�c����[�h�Bc��e5D�	�8�FT�IRX�H%��(�<�q��:u>�Pĉ��H���ȟ���ݟ���Xyr,�q��"S�'�<���G�}x��Bk�`[6�j�'G�6m�O,i������O,xlڶ�Ms��K�g���q��'GAi�m97MP�c� FK%d���-��<Qc�R�h���]	�=s11O�0A����l̲��[Y����#YD�̊D�7P�9 %o�O����OB�ɓl�����.�I!|=�C�T��03Q�����Ol�D˧u����"�<I@�i[�)̊�y"홰/*� ��B�G*�RD���՜E��'"����R��|��A >�u�牽j&p����3^����
rE�0��l(g�^h�h1�U ',�I��?�&�Z�T�y@��?q��X��ȱ+X*sفP%�& �H`H��?a-Ox�aCR�NH.ʓ�?Y�'��SS���3�Y���	�EX�(�7�w~Ҭ�>��i��7�́3��	�(B�Hx�Ox�U3�ڭ.�x��@H�C�J`+�G��1��!C∇J��Yʛ��L��y'B���d�$`��	�7-�89v�ÙaŠ���#m���Ir��˟��i>�	џ��'��(1gg��A���kZ	�b�#b 9e�a�ע�jy�}���d^*ni��=��Du�"q2$�و|�H��@ , *��$�Ͷ�Hv�ÊBd�ɰ���3����2�yR��3�b	�g��%G�"QR�o�.�?�$�'�Xy�tJ��~���'���O���Q[>I��f~�2%��L p+ʅ;�0��t#�ҟ�����`��-���ʟ�k����r/B��́#��8�*�F�i��V*b�� c1�O"���&�<����
���]�n��p�rg��W��铭��쭰SG��<Q�C^.1�T��ߙ;t�p�'F��䀁F���"�O8���M���i�-Q�ku��i&��O��D�OF�D�<��A��/������?�����\�dܬk��H;�eݰ����'����~�d��unz��C�O��rg�-k�ء�W`ׂcР@b����$H�}�1�'I<@:fhۦZr�@ %�J�y´�pd���'rM��܀�P[�E'�J0C�Aњo������,��?d�� ��CK�S����I��`�,H�P� ��[�Yl�`6k���� lݢ��'�<7�O�Yy����9���Q%��	g�*u"�<&�cB㜭G�����4U�BQQFH�"�uG��i���7T�=Xw6UY�ˎ�
/x	��n
[��be�\u]���'�,�dH	A2ֵQ�I�O
�$�O*����J0L�T�Ω+֬ۇ��u�:=`QΤ<��+�0�l�����?���"�iD����p��}ң�;��@�؀b�p��'&�6K��5@���̱� ����6�������{�d�zD�
���S�[��ts �}��b�G6?2��	�Q'�˓:�B�-.(�]9�Afl�J"/�=�L�q� ^��'���'(�S��Sw�Gւ��ʟXku�1O�V��!N5�J��& ���ܴ�?��Z~�̳<Q���M��*�9C#FQ�$�yV�Xq1#S�>���T����H�`���<��B\�O H��1Wnr)i@V>y �;txhx����I��qA4	�;b�ށ��)A\Lh��?�����`B���缓4�Dh�E�Y9j�) �(�<Y��?y7��0ʔ��'m�6�O~ 3O�{�N�G@�h�-J
/���f;;9���!KӪ	#��v���il>֝
U�.e�B�6��gj���9 ��E�e�9��Lj���Z����'߬��='��h���O6��O,ٺg`_�#.���Eϰ#�4h��m�Oz�D�<1����i̓�?������Ef�M��lP7��t�VB�"l�.`�',�,����l�05s��OV�Sw ������v�0GŐD&�`��[kn:`a�H��`���Q�y�'i�V���v�j�j,OZ@A���b�H��ƄF��9�3�ӟ�I%�\���	П�S̟ �	By�f� ľ@��
�pfR9h3��Щ'� :{B�'�L6M�O$L릞�<r�O�Ao�"�pqeJH_����!��d:�4*��8�S��s�>�KO�<���̃%�R�:���ڳ5O� i��@�+��ڣ�ٳ�hA��'�
��D-��P���O����OX��ڍ:���'qC��J C)ʒ�sDaͱ(�����:(�а����?�����w$��|Z��3���w�*�aׂZt��c�Р�-���bӌ�n�����(�D�谞?�#/�ֺ��M�m� #E�>T ����`��\S�'WB0����Pp���ҟ��"f�=T�jU���@��� "4�n�����2}Bʑ��֟��ɟ�'fH8B)#+%R�'��$S�X蒱+�Of�,!kҁ	"L��*��dQ}��lӺEn�J�$��2���f͐E�N)��+��d��$���t�dܒ4����F�qY�<��3O���N@~�D� �TH���ΔM���r2BبNZ�L!&��0�?���?�e�-l8���K~���?��Bu���@�6�1�,@�+�<A��^���5�L6��DVߦy��y:�Ӽ����!^���$�<)��@k�d�˕��RM�a��O���P��D��.�������Ӷ$
�N��)"#�%4 ;�,��I�8� O�+����됀F<>b\Q�I՟����?]�#i�4$p���%����P��Bԕ'��+���y"�' B�Oe��O>�0D� $t1�T*\d -�D/�O}�s�
�n�&E�`�	!E��$���^����i��Ң ۩ 5V�R!���CH����Į*��X 07O���kA��?Ѣ,G剐�?y�0b��xv�ӓq*�KCBJP�B�*bŁ��?���?i��?Q/O��t����DY5$�QpC�>����	�����F٦���51�.� m��=�MCG�i��܈E��82I
���*
�൐�h
CSH���N� �'���9���޺+qa�ʧ<�Gg�qR��aM G`��#+��E�|��A562�'���OW|�֕��wܖL��0 �� Ď��/��j�'P��'�n��3K����ĆҦA�	8'2�W2 "D,J+p�(�zq	��k�$i�g����K��2�jYoZ�?�B����#3�T�f�R$� /�E#��K)bWc�H%�e \����e������c��X���	ڟ���"{��e�㬃���9��r�������'Cne!գR�y��'h��O�J��k7�@�Y����.I���'cݗ��DS}"}ӾmڨT��	�JuF������0p
U�ܫF�0����
,�p��eJ�z4D��I���x�$9O�֝�P�m��[���,Oj�ˇ�C.G�TZ fC�X�r��C��H�f啳c�P����SޟT�	{y�Lՙn�ҭ��i��:�,��@nɲ ��E����a�剷�M��(�08�'���?��O�Li8��d�.+�:$�a��?�f��/V�qk��G���͓O-F�0��~݁)�f:fX��?n�jL10E�('π��bΆ1k"C�OȨ�r&��nV���O�����2��2ɫ|!郖j�.��%�J�+"��w�������A��?���?I��p.��-Oæ�!@�r-pq�<Fe���B��	S{�����c4㼟��,�U���!�\h�;FsY��Gَ�R�ӯC
��B�ԓ�y�m��j�8��	,���q*OT���*��:�[ޟ��â�(]D��J�1a*�5$�ǟ������Py�,]� ��q�ET�L���+�&�;t��<v�!�T��{Xm��l���W������	�Nʦ�� +���ބx5�yS��+�Ѡ3�'������x�o?���P>)xwC�O�L��!Ol��q��őb
��V��)
H����?���#x��;�Ǌ���'�?����?)r���g�e�q" 2YNp��t�[��?�g$E	
j-�-O�<m���4jW�9?�;H��qY��V�2S�lɡ4��Ђ�
���h�i�B���`���Z�t��)����KU��n���Ù�"������gX�`�,Ot���&1-fd��nO�V~���򟀐�@(�<n���Lxm�v�B���B�� ���?	���?���]�`�(O��Yƭ��{�ԭUL&tˊ���$_}�DeӀanZ�7��	��Ea�?=b�Μ�>툥;Q��4T�Ĭ	!FX�F����s.οZ��牛�zhpT�'�h���<��'r���b��t�xq�"� *�p9`�`��Y��'��'b�'��	�uM� ��n�@��B*m%�ubˤ�Px�è`�X��4�?��E�C~J�>��i�6mK%�(ȣ�&`< *V���ii�d�87n�sq W|��d[�H�,�[w�B0k�!�}�d����5{Q�M-@e! Ƭ�y�
5���cG܈���O����O�����p����Q5YW�QT,�r�̩�P�K�P�˓�?ᖏ-zZ�M�OO6M�O�x38O&���O����*K7?u@����Z����:;i��b ���4�L�f��N"x���I$@�I��`������	X3B����Siy��R�	y�fFbm�r���y��'�2�'��(2�a �b�!n�� y�'�"Z��/����I韌�	�?Ͳ��ܧ!�����h�[�J�"B�Sc�(��	5�M�!�i*����'=a[�N��|R�hð{�(�I�)ݙ%s*�y����{�+ݝ]�����d��<����$�%*�F��'�ĴZ6-�&}���2e�4+�q�U��O0�変<���D�O��O��d�<���&6f�3�J,�깱�k�� >x�Ra]m~��v���A$2�ɟ��DjӐ�R�iZ�$ʽX�������a���">=��"���6L����7=� s1���ؙ�U<�y����-�z!��� u���Ƒ�?!E�'����G�U�?���'���O`|H�Y>�K3"�rcNy��I	��5H��3� $���l���	����S)Qp����wR���^�̒��n���&e��$o08���u:Q���?��qe�ԺCq��%��ܚe�Ӄ#�
Q�F�T��Q �'��l�Սǟ̈^'��#�B�<6�����'�iY�[9x�v!`��<c*��(!�'H��'BS��Y�� �K�P9�I͟��ɼ3�-aR�֨@���Ai//��IZ���EV�I��M��i%r Y�'Z9@�yW&L+7'�&0d	�v%���ޑ�q?�ir�D�@W0�#Cd�D��.�?	����M���2 �,���t��F��!8�O�O����O
��׏] �Z��J�d�O���k|}["H�lо�8fΘ�s�b�$�e�uc⌻<Y��i�R����4���E{������*R���X�y���Je�[���Z�[�/Q*I�;N��'�Υ��κK�.� ��9š4-T��E�'��XA򪁙yJ�ɢ�?AgΛ�*H����?���p�)G���� *s>5J˅]^��,O�X%��F�>�$�O(�d�$9c��<��Y&Y�}��H�q�@�sO.+7�	�M!�ix��Q�'鰕;�^�$�� k�HyA�+ː1�:��s�R�1"�4
��ԑ>y
8��'�\T��O��x��� ���Dϟ���F�1_�@����`��0�#�"0�P�R�XП��������\�'�^D�k�~�BI�^ u�'��7^��Ջ�!�yBs����5U������������4H{��X�/E=\LcM�}�d�HV�4P�qH�D�d�̓R����/d����L
)P哧�����Н9�ʨ��Z����/�--���s-Ȭ�?Y���?Q�'nT0K~λ~�^�Q����H�BQ�v���wr,����?���td�t��k���������I
N����5���g-[�xU���V�ۼx�.���$������L��oz>y�]�� B-d(ϓ�Y�%�!Q����`�(ZV�Z���T���ϣTZE�'�X�dџE�4\�&l�O��d�O|34��{'*��n�� ��13��O��d�<���@� R*O���ڸ����8֎@��N%��=��	Z9Wa�	9�����5Iڴ!Ѿ]��E�έ)|�钯&�r2b/ ;g\@��ap&A��I�a���� 1Y���Oc Q��PA�O8���(gP.£I�E����˟�@�Q�U
�������Ο ��Hy%�+dC Р���"�b��0Et�k�K�^�I�MC�����'_��X��f����J<�B�9�tIf���7A�7�G�&��"1|��D��O���M��u��λH�B��D�ư�@I�'t��؀F»O��e�Ʉ�?yA�V7t�����?�������L1���Q�@�R�٥$�18���R�$/kf9K�bF:V��$�O���\��"�<����yw�� r��E򃯁4.k�#Q��\GL6m����c ��\���J�0�B�I���i#r&s�!)�AE�^"�4��+9�ԃ��~[X��B�D�#�O�t�ǭ�vy�
�O�p&�_�TF�����=$�S��8� tꟕ=���$�O����Or˓R|��-�?����?	�@�Ύ�Ф�4b1�@��D�?�2�KD~⍲>��i��7�=���DI�@يs� :����e�;|<+H���^�v�;��Ƕ�F �'��N� ]��¡ _l�`�	L6*ѲA� &; �؟8�I����!���$$?!��ޟ�]�G8��	)5� �u�K�.(�	�5�������ay��f�������iޝ#�g��v r��lOI��<)�G�9Y�H��2Ł�M��I�8�5�]w�8@a5>O��Ċ	�uGʎ�U��Y���`�D�i�$�L�� SU��^y�i�O��[�o�	e�d�OB�D���i��ˌ�L6`t����j��x�&�v%�ʓeE����
֙�?q���?���wKz5�O���%�̮
�xd4HϜW��`��>��iC�6�>��䜃<pA�̟���t�@�\}�i�`�t�=��n�+#k���<��D��b�
��\�5�2Z����$lhm�d�ƯUe�= ��"Q.�Uk�ɖj��dH���?Y��?�����Z�i�:ᓦ��O>4A7k��$�mܲ�
G5OjQo�ݟL�n7?�]� �	�]xTG�(X���rϗm�VP��	S�|4��II�{�z���v�������Y����r&xa�/����8l<��ۄD��pځ �B��N�z���� ���	ß�	�?��N�x�s޵���;N�����Z� CP��۟��	��48g�E�n�n���$��4�?9A$�<�e�$C�6(AE #V4���j�%[Ru���	�銵�M�'.[Zw|Z̀�2O��5��s�^��ք��}����B����L�mXz�ɑQ����I�����T��?1��?!�4 V�\��0B	��g^8h��'>�	P�hp8���ǟ���Ɵ��S�j*Α�di�!)��ځ�^��uڧho�	���^��ܴGPTM���8"qj>��lɕۂX��_0T6�\�¨�	7U��"CO�}��.n���O�f���gHM�u_�,	���4פpic��p�&�)�?Q��[\v4����?�'�?i����As�yJ&*�[��q�_K���xWh�&7:�I�*O�hnZ���H�;?�#Y��[�4Eu��ZRL�%oHT��F'[�5�dQr�iC��XǃP�(@�G*Ʈ�yb$X�uǖ��;
Z����%v����פ�$���I�q茽��C�O�T���+Y8-k��8�	�x��
]��O���Z�
�h�܈��X/{M��`S,B�c�HRG�'�b�'�������T�'{�6=�|!pMˇb?*����i.��`Hז4tlZ�t���
 ���!'�?��ʺ���ݢ
(���4HKPQ�@��-��E�'�V,yce���P G��%���ԟ�zr,V�VO���	0EKeBG/̠1�,��a�Z0��e�I�h����Е'�v5�p��<��I��8*ub�bF����*D������D���!?A�S�ă�4Aכ�*��~2hɇGb2��w�I��P��`͉z�.��Sd�<����Q�]��o :E�j��O+|�K���� ����J�t��d�5!�T	�X�a����O��$[#(�ǉ$�i�O��D�O( ����,d��:� �V�!����O�T��N_�W�ʓ���'�*}��O�J5�<X�A�:t�(㧌�
_�� el^�*�o�!�rpKe��̺�mA�'�����gYĺo��"	���EK�Jk�Z��� $Btxap�My��O�I���u���O��D�n$0ǉ��W���2e�/9^�kAM�+�6˓�Ps��+�?���?���t���'�?!u
�Y���3)Ŕ~st��睶��$�O�6-f��2CV+'[��
��jI�iXw�O�)(��lJ��D6�M���
��yҭӝ..��̓~�� -OD��	�U�����/p�,�f��bW�aĚ����O��d�O����O$ʓ7�Ա0����?AQ
�	Xʼ�n�/q��s�hT��?y���?��K��<I�����9{�4��]9U�ݭ9���7��:��㷀ʬ >�{���z�d�شz����ܺ[盦)�hWBu�1�;E�X���̶��UjĀ��B�Ȣ�4�.q���?����Zs�S%���k�i�9�tV�{��J�������O��cbL�)*(�S��M[�WKhΓq�dd8p&�f�I��Y�
�]:�	�H?	�M�+�$T�i>QQ����G���yN���� T��A��o�TC`F�q`�i�S'�!�?)a�1Jn�"�?�C��#? حX���?9��D>���q�
S"�,����x��݉���?�-O�JE��BOJ���Oj�D��:���GE
�����:��1K�
Oe�� ���O�_�Z������tҝO�؈@��v�z�sF��� \�'����0��W�W?pC����rg.�ٟ��!$�����D��1�^^�=�3e�"j7���'LQyq�^�y���T�'^�T�$��K(�ly�#��<M�1�4l#*���S4wybks��D�<�	���D�O����a�
�� p����G�O@Jɜ�s�&�&bG>w���<�"�9^w�ɱ����<��1,�5CA�N�Wp�}�@e�ǟd*�E�Lpu���?����?��'Z=`�H(����ǂC�Mc6�Dΰ3��M�T,�:Ƥ�O��d�O��	K�˓(䛞w2x�����)�ja�ئ�`D� �'�2��!�~R��6n���O]H���ą� &v�ٶ��7�x���b�>�Q��P( �'6�uE��<�5�'�а�¥�l-ϋ�f�,����5u��(W���t���'W��'��ɼ")H�(�J�۟�����@"��Y�Xj�̏XA�8QF �柼�$)?�#\�<��ȟ�Eŵ��X�/'^8��������7J��+��8�y�V�RV9{r��=�nɑ)����'�*5����O�������)hl����
.w��T��ߟ��	(�l�r�o�D����	ß�2F_�u,�=�Ql�D�\��U&�͟L����CD�1�'�6��O�P{唟��F%�P
���,��Fb?�^PBu�W�"�B���0k��a����S�fL*�yl�;;h����F/��EH�����fۛ@�����a�~�m��L���Li��'�r�'���H׮p0��c�jI�&&�� !)�� fW�h V.�1���Iݟ��I�?���G#?QŌĢ ���	�R�0�"�R/N��	��M+����8�~� ۥT*��Om|,RR���D	tm YB�힨Z�N�n��y���0�����*�BD`)O���ɀ�L�� �({�| �u(��Q��%��oi/�1�Iӟ��	ӟ��	cy� ^"?�`��'p�8/�Ҕ�E�	X�;��&�y2Ap���dătG�I	���O�6mb#h �2�K�f�@Q��%�w6�T�bNW�?X���CL�y�K�2$�Zw6Ua�����P�Q�^�(b�9�(�=��T"�m$V��Ypg��OX���O��I6}�����7�@P��)FT�a��3���O����yX�!����Ds۴�?1W�@�<i�x4P���?-BuQ�&��D��v̉���Mϧ'�ȡh_wFQ�d2OT<cQ`��x� �S��[�t,(�L, �XH���bڸ�ڳ[� p�OyP��vL���?����?9���+yƬZ�#�5NpI��E�?�����J�9�X�ʱ6O��$�O����<��a0��I(��y�խ잁@p����O�l��M3g��A?��ߚb�%���f��f9Q<Bw�:�`�&J�|i��'VŔ�	ߺc&"ßDq�Iʚ��d�6¼Q�R�4|0���sg`��/9o�qh�ӟ��i>���͟�'b~�4�2�|��d�	;1�|���(�b��(�b�'d��f����S��#���Ц��6,�f�̡4���;�6�)#lN��M�pBԖO�\`�Ti�+K��Γ�tii�}�UR�#��4���N�@F�t��k	-���Q�mQ��K�Od��MOt�6���O��쟔��'�|���@쨼�$k��
��H7W`�ӓo��t��q��������?u��h>����M�;k�r�ڃIJ"Y������$(�N��r�i�67M�����&4��P͟�l�Ҋd�eٰ��4�A��j^�FJUPq����|u͓��-���O�a�S+EyBg�O�@��0;lf�]Pݸ= �U�N�6�1IԾnf�d�O����O�˓g\00���P��?����?�U�T3���y0C^;(6�U�"���?Ya��O~bF�>Y"�ion6Kh����#e:��h�A(]��D�7i�d�$ɱ7�����t 2�ap�ڡ �'[��)��%L�uq���Uhȣk���ƈ� ~��a��T�	ǟ��k��	<��'?m�	ϟ���2c�Fy��+�(bdk1��2و��	g%���׌�����I?�M��|Qt�yWg�Tiji�C�P;OJ����ԃujh��+R7펩uJ���g`�e�&���<���`��ݶ.���A`kJ��e&7�D`Qh�d�I&�?1��A�X���?���beG�Z��0�S_+U��eI;֠`R/O,I1���N[���O�����0��E<����U�v<���#��V `��E+�-�4��'�¾i�6܊�'�V(ʶ�e��'�7<�<u�#��K�~Ql$Q�Rm ��13$"�q�'!⢨�ştCTF�'��d�㟼h��	����`C�� �.�JSd�²�ec�̟����X�	˟��'�t@j���_/��Ǭ'�\��/W/}�H2�N���yBmk�����X����������!��4#=����A�L�C3�S0R���q�Ùn༝�Wa�E�l�s��p3
�A��c�U��߾n*��|�a��;xP0@��S�<���$4Q$����D�D���?������͗����S5��{�e�q �+3*X��F�F�<���?���)j�:u�'6M�O�iiU<O�*$nծp����ቊ�%����L�(��$�%�|�Q�x�|����� ֝�rn�]x�?���┽.�\��C �K��QY$j�q��'!>��3/�<Q��'��x:��ץA���'w�.|T$�ȴGY$r��I�Q��_���'_�I6{g����}�l�	矴���&�0�K�	�SP`][����Y�Fp)��4?	7X��;�4)+���!f��Vn-8��O����iE���p�qHL�3oHuԌ��`�Ƹ2Ү�/��'���G21���j{h�`��s$�&=� at	[ �x�i��'��h
`���R���t�'=�X�`���&v �.1H5|3b�+z(�ԸE�??��i�"	χ���X}"moӈ���AXC�cb5(��k'� ٦%c�b�#5J����j !g�扳d|T�F�����wD���y"���2ȋ�W -�l(��Y6�?)��'���B��m6�'�"�O0
�B�P>%"��H��M�M�zՒ�V��h�Ebv���	� ������AZ��w�H�q���<C���ck؀`�%:0�dӔC��m��'y� �a,�`����h����0o�� ��9�i
 L�̺��G�j�@��7O�̒#K���?ц*T�
�I��?Y0o�P~:�J���"u��/k�°�s�%3�,؉��?����?)OpQ1�/B4�ʓ�?9��J�#4����=v0*# ���?���@f~2E�>���i46M�z�$�$ɼ5r��x|JX"E,��S��� ���y�G��R+�M���ىo���j(������'>�գ�H�<C���@�x|#6ȃ�zM�I�4�	:g�
���Ym��<�i�т�L/�IS��<��ъ��6Hv�Bt[-Oao��xb��1?�;B����3*צ�������dΌ�"�R3JD��ZB�i�0���#�(K��N�6��I�xqz]S�����w�&d4`F�˸�0 RUI�<HV��0/O�����V\�TmHџ��	��L������	�ኩ1�V(�����DF�qQ�Oyb�P4t]�Yp��'9��'����P�����'�@)c�٤R86\(�Ĉt���XC�>��i�6mW���dR86�@yִ̟�e!�7cT��n߽K ��qM�?c}�6A_��$@�)ّ�c�vm
�Q�Xc�($dDj2��*X0�-���o޴��-�6�rx���?����?i����dX�:���"���Ox�@[$�J����jG`$(E��O�en�ȟ(K2�#?�Y�4�Iæ9���ͺ	ͺ�����n�8�hF(9�1)�lVu���0o�ڟx+6�P���N2���y�'�����)sd���D	�AjO�Tک�F��8n�yJv���H�I͟0�S�U��X'?�]9hjY��AͶI?<� bK��#3z��I��\�	���A��O_yy�ns� �d�>	��P�/g�"��8}�D���iuy�U�O�S�O�/M�6=�b��sݱk����<t�{�pI���e�H���<#�ڽ`'��OB�PD�Ny�OH���o/B�0���O��䇍؁�To�}؄�0v�D�\p����O��"`H2��$�?Y��?�'%(�h��G�V��V��A�񢉔BE������Ԧ��ܴT�vq�%�8��w>)�""ُm������+f/�񆙳 ���
�f�1h�b�Ag���.Pd���
Q�<ʓd8�Հ�l�&E ���S�ژZ:
M�U�'E���-`9���D�' �R�hU�Z�`Hy��@�w��b�/S�EE�����"�M���UTZy�'���U����[rŞ�+�~�Z�CާcNB6- l������P��L�:Oh�R�I��uwlU�$x4Y̓|q�2��Y1���X�'���>��I�?�a%�5������?q���"��@	���A_h����8=��b��0.�}"TnT$�d�O:����L ���<���yaU��ZŉҬ�m��%�"�R7���;�E��\'琌BZ��;]R�Y�;w��L��+��\�'��(E�u�\.�y�k�������AИx(O�-�	�)ʎ��jF��*`)Y�_)Y��� kI�̪���$������iyR�]�}z�r�'���'M���c�>���%�2�XUA��'���O>��'w7����d��4��m��h�����O�4)��)i�!f��B�7O��H�)�M�:�J������78�d�%6�`�c)�6�䥊E'�!=�Zݒ�	_��?����?��j;o��9K~
��?��1YTU��x���ֵ	�(EI�oX���١�?��*Q���'�t��O��,Zc���w�;vt��p�'}D�\Чk�\H�o�eѺeY��ݤFi�͓8~d�J�����N�(�zi�G�Q���9"ܫ<v�Y�\��i�>�^%�Q[�?Y��?����P��!�� nGX ��e�Y 0�IG@`q�'o�`B�H�)���'�R�O7v���^��〩4>r�B��J�,����ǟ2��$Oڦu�ڴ�x���R�~��W�$�w�BRȼ��&�`Țӆ�(�� ō) �l�;�qɁn�O�|���Oy2��O�E��׺Br���i_pHBx�(>eG6���k�O��D�O���O6����@N��?�d���[�8{��˥&��?��i�r����$@~}r�f�r�m'b�f�a�G�, uJ4��a��UC7;�v4h���oVh�	4zp�����q�+�#�����}Ӣ(�"��t��}����D
D:	i>�ɕ/����럘�� ��&?睄��Y0�ϐA��d���,�E��ğ4�ɋw{�����DyGq�J�� �^��$�	Nq�ъ`��u\h 8k�*E�����OJ�[�oM�c�P7=�n/�2��S���n�I�cѓ�0�y���
d�O�*<�D-w�d�'����
�u�a���?A���?��f�4k��I�.S	��9�"A�?�����d���d,ʳJ�O�D�OB�	���ySԆf��)&��.3fL��S����O��nZ!�Mc1!HC?!��˹]*
��l3��v(ʢ1}����oJ�ECA@���DC&Ƣn����l�a�'}R)�A�<I�N�[�f���FGh\N�*��I�/!0���'��O���'�	�H՚��Wȝ˞!��ǭ\�Lt�+��5��4�ݴ�?�2�V~�+�>��i6��u/�$j�A1㚣{f��fm{��)x!��Dp}*$�Caf��{��[w�8m�5)�<�`�`�"N#�fe	P*Ggi������@��Ԑ$�	�0�	�?Q��K�D�Ћ`0�t�
��z���'G�:(���"`����'~��O�x�i�O�BDq��66~�д ݉�mSԠDC�q��Ϧ�#1(֮�8T�������Cr!u��䣁>%���w�U�K��#=��}ϓxj�`��Or)h#o�|y,�O��kE��>{���)#���dKT���s�ΞZ|����O��d�O�ʓH�*)0���.�?���?�@����s3�,#A��r
���?QbeXD~��>QP�i.�7͉�C��������V7!�H�i�/�h�@��%Ф�.yj�0!RE3���mZ0��%�^�<9[w/z,���@c���&H�r�u��Ln������M	P�>��OV��׃uDFP�0`/���O����OAW⚧���� ��@�d�%��O�5+0��	p4ʓK���'_,EX�O�nٵ=��4��Y3%�rY��^�C��
U�X���%o�J��X��FѺ+c%H�h�bD >��-��kb�m��Hߕ^��<@���"���3��&;6�yZ�l <���`��'�R�'Y�DM��,wHՀs#�u_�����4:(�aWU��y�(�&��Iԟ��I�?�WO�Ny@��|&�	R��\sP���#ŗk7$�?���n��%�O^�P&����ɜ�� D����L�"M�5���JIX��A�
�<��3O� 2w��?���K�y)�	�?��V��a@t!4I��kȧ((�`�q�?a���?y���?�-OR���ݿq���B=jξ����MP(x�BQ�m�\����I�|���i��I��MCv�i�Ep�Bq���y�I�Y���{��Ą+/60@�Y72��ј'y�����Bۺk���'���'T��o[�-��7O¬�yR�C����權0���'�2�O��$`���w�h�'�L�
t�:�)�6��ݢ�Y�`��)y֤tⶭ4!�i���y2� ?�%j��ǖ#D0��]{'����'�� y�H����O8�5��[H���''8��1y�&qs��=>j�; ��F`���'�>U �î<���'�n��B�P6k�B�'*2�]�U!�Ѣ��{Ԟ�j���l�r�'�I%G�pq�/Lş�	����S�,hm*���%K�v�q1FM�v�1��;?�bR�� ߴmG�6� �~B��&��	Χn��l`b�"iB��
�2N��#�&TW�!��h4��?��e��OBٳ �Qy�����!�$�A0d�j�h��.D���8 -~��V�Ob�4�����Oʓ@��	p�m��!<�|���`���mY'P[�T	*O�]l矤
@';?a�Q�l�zk؄C�ƽ�vM��`"����4�0�b ��?3�[%k���?)`�T-0=���l�P�?O�Q9'��6�d���߇-�,H���'��D�~��**�O��d�O��	Z�eh�'t�f�nΆiX�b���Zқ@�P(`�~u��'	��'��\����.Oiob�e
&�˶f��m�Ǌ��F�P��@,G��M��i����'�d cŃ�<���'z��8Yw�D�Z�ϒ�V�"P�hI�h.a��%�X��R;Kw�p����z_� ���<�p�	��+�?yT��!I����DԀ)d��BFA��?���?y���S(y99���O���O�3��"��@���č	,�:�L�O���ҕ��R�OܵnZ:�McQ�[?�DN�=��p�Cv-`!��J�z ��k�p�bK �)�dD����U<˧~נ �I�fM>��v�4E4 eq�K�d��,�(,F�'�\��Uz%��T�'�2�'f��zc��(�����8
"((��'K�e��	�MS�u2��ywlE ���!bi@�	���r��Ǡ(:�$X8,�6MݝS4̤
�&j�;¦��<yǍoC��݊�x�q'X/L8�X:E@�!m�4��לy���>�?a�� ^������?����bT�( n�p�oUR�t%ʇ�O�N�ݲ*O0�� D���lʓ�?y�'*>��O0��#Bه��ICG�G%$J�hb`�>"�i�~6�ũ#����8Ov��̟�̣ EYC�b���a��Ru��D��aT����d\���p�C?�99�T���S]�������l�
@����: 6���a��aA�H���?���?������?����d%�OD�IWŖ4b�$pJn�{1X ӆ>OioZƟ���=?�%]���4V���������1H��\����c�9s����v΃�0F�Z�"R��yhD�m��௻Q�B�3�ļ|"��w���� �[x	B�"D�iަ����B!j��'r�'���@�~#��y��٥ ����㋻O'�|�BԆe��'<��h�~���]��ڴ�?��d	�<�r�O�J�r�pG���8g���-60��	�\рOE �M�'
\��\w���rR7O�����= ���	̤\�B�(���C��bX�U��A��+�l��a	څ�?���?��'�D�r�߽$��/�?�����6]lՙ�!�O����OJ��V�=vJ�����,Fxja � '�|z��(O�dl�h��e�Ord ��E�����z;ąTmӁ�
�j�)F��Ѩw�ZO6y����y��� ��Ɂfj�L�)O��T�<*|�]���Fy��f!�ПXO�8��E��ȟ��П\�	Qy�$Z�% j��1��$`��E,/Ͼ@a��* ��'B@6-�O�� f���A)O`6���|�7o��l@�n��Jyn��V�;�^+uAz9��la��h @E1=�N�<�� q�'df�'�0��pa��GJ��ݡ�����7-�����'rB�'����L���	þ0Iv'�6AGr�y�Q	�r�	B�NU�e��ܟ��	�?�K(�vy2c���{�x���(L>��Jc�ċ8	��l���M�JUR?���ˑ,\*�'��P�]w�JdjDf�2���w!P��d�V7-��0t�4�?Ѥ��0�剅�?��߾z��h;��^�^h��G?x.��p�	�:��Q���?9��?�(O����X����OL��V;0��@ �}+J�Ѡ�0�`�dޟbF�ɚ��d
ߦEݴVǴi���@�ig�V�*A����E�b;�@��h)R�ɋ	@R�q��C_9Ι� ��|�fF����xu�-|�]F9W(�4�`h8��m��'b��'Q+���^�OG��'�"��<x�iJ134�T8�͇J"R�|I�a҃�?����F�'�h�O�A7����p	D�P�9)���t��з��2n�(oZ�&�́!d��sb�\��yb�ڶspv���n9.�:#핛
��pp�dV;���a¬�:FD��&^2j�k��Q��'(��'I���L2�R睱@hX����\����SP�P�s,'w����������?�9�Lzy"Gֲ*J�u����+jE2��ȧ$Dt��?Y�WE�t��
@tI�&:2�	,�Tp� Fڛ2��Y��@	3^$�8�q�@͓d��h����OT�W�QiyRB�O�@��N���@���%rw�H�� ���pAv��Op���Oj��O�ʓ,�"]r���+�?��AE~�Q�#��3@�5W�\�<�`�i�Ro^��D�_}R-~Ӏ]l�$���Q��R��=Ӓ��c;�ɨ���\{�x��`�sk,才1�ܑYG���`0�+���)��ɀ&�җN�P�g`�S߄��lW (�y�rlL˟��I㟬��ma45$?�84(*�P6��9 h����^:7?����ȟ���?j��0өs>��	4�M���$��	Pm3�d����`R:G�t!��a�@?iR*V�fPL�x�4��.�u7���v���䂋����)�O��EZ�+X�h�L�KP���?��a�M��?��f
-y� ���?��Oo$Tc�ėW��,�N�38��h��?�/O(�!�3����O>�D�.�*��S�|��Eؕ��<r��qK�d,�I���D�ͦy�4zd(��XԠ �w>� ֌z�� `��a��}�Ƙs�ʍ�n��(�vGb���#ah����e����P��˓`�b����[�_��@��[��i��'	(��bO�t2�����'�bR���%�
jeb `X7p� �!�͓+�&]���S�|���M;�"Hl�'y��M{�`��4a��ϼ!�t�Bکw�f�\;b���Ș,�u��'R�0A�޺oڰ'�m�P�pd1�n�?h�P����n�
�����?�L�.%�L��?����mՉ��ɇ�¸�֭�3{��`B�Z�4z"��Z����O���jq;e:���ަ�]iNVu�0@_�[�hu3t�0�u�B��M�ұi�l���'Q,�h &�f�Dg�'1�Μ-B���+��;"�"�WA�_Âl�R
���u��p�d��t�˓5�Z��kR�'}<}��Ă�>�
Y����T�r�@��'T��'��[��)rE������ɼB�R I�+�0/����Dz���ɩL��"���	�M� �i ��8�';nS1��@=jc̗�K�,� M h*�4����"�Mk�"����)@���$jR��� f���Ӧ1�:�)�����D��ݟ�J���ˠ�&?��Iݟ�]=�VH�GT�]
��v띁%����	*VI���4�ʟ���Bb����1?ͻh�&]�`O�f%~�Q�!�	6~H���Ds6T`v�i�>����ڝ2w�T#p�	#F�f)����&N�&B���2A^g����DO�=c�}{�_����"��M���W�?��?Y�'g�X+��Mgta@BF�_�f,�5����!BC��Oh�D�O��I��i^|�}Pȉ��ڼcY�Dɕ(�r��I`�U��ڴ<��n���~��A�m�=�Ot� ƅZ�e��ꓽ��ĩޅF@Y�G-��	���K����d�Oz,c�ǐVyra�O�x��a�Ds�U�WAڸ3@șį�%+�RAK3��O����O��d�O��yuҨ3̟�<����8�Xe`灂�s����a��<q��i�be���h}bK�8tlZ�U���؄F�hī��ǋ��y�S�lil�z�ͦCaX�I6D�2�҅��޼ˣ'�o�t��ƭH�ڵ-�f�@�C��+��t8�Ӣ;��0�@�O����O��	_�m�V���.T ]��f"�"d$ڬ��G��d����O0�d
n��]� ���ܴ�?YQ ��<ɒ��;q"�E�խ���f@I�JL )�����(�D��$l7�M�'iǼ��Xw�^�C,�O�0��Ey�ĩ��fǫ\�J5	sM}����<�t�SW���0Ξ���I�?)���?�p� )r%�4qD��;w�2�b���?i����!�9�8O2���O���� /�}[b��YKZ�q�������Du}��toZ5����b�(������F-H�F	��A����֐E�N��q,��LJ��"�<On�݊al�Ē;iy�(�'� �[`JЬ���D���|��� �>O���3m_�>xaz�BVm����gL��5yJ�+ț=~?Q�W�y���'��7m�OJy����$�O�}l�K`^U;���j Ɣ!�'�:z��)��4t殉`��g�>P��\'�?����-�H�}�hd�Fg����	�brsʇr�	R�M�Ob��	/m�� ��`�I˟��Sa���O �3��������O_4N� b��j����q�'>��'�TB^�O�剀�Mϻ]w�˴�\=X��С
��.�|9����?��`?�!h�G���lX�:_w��L���#�Ba�� ��!,�Xz e+t�d�	r�J�0��z\�WU�( ��r�-X�$��<I�GX)OA��b��|�t|��D�S��"2�۹�����ܟ����;�<�aed�nj��vD�"������9oz�^ �Iܟ|oZ�k�6�ɜW�����:�>a��H>Wܘ,i@�S�AO��$��L0����,�R��5O�ם�}�����@$H����ձ|��A@t"���Py�@�?���?�BgV1eOp�K~���?ͻ,TI�r遭�t%��/�/+�:����4Č�s0�]*�?��$�V�'��`x�'T�w���>I
��`�X����7-~��s�D�k3�]lZ�V�r��S�2c��bX@ٮ᯻H>��:��g�`�0!
&`��?C���fV��X�/a8� ���?I��?���dG����	I�t�t�ò�d��Q'����(h�Lk&��O�D�O&�	����)�OR\�B�+�j}8�
�	5���!t��G}R�c�0�lژ5FJ�I�)T�Bb�`��\)< ���g��3�xe�2i��hjg�u�X�	���X���ݖM��$�	M�z�X�DL� 4��0�ӓO�p�������bA;>���'z��' �\�i`O ]��I�K��A�HT;=ư��Bٺ��4��?�M���`+*I��?�F]��Qٴ%�V�REŲH�����[��J7DX��A4��(zϬ cD�� *DܰX����J����<AXww��Nltά�ӆ��i;J�ڱA�q�53�� Ո���OD�d����
��9�9�n����B]�q��6=:�����O(���OZ!���D�p��O�!mZ蟀��Ej��G���}��C�x�R<I��~���	�r�e�Ƅ���E�Ӈ�
ծ;�����'G"�#���8�$��wā�%4��k�ƻ-�h�	*`
�YB.OH��	g9t,@�ǟ@�I�6�r�C�H�h���4��&i���<�'X��VA�(v���'��O�VL;3�$� e�PB��@^0$j�ϋ�y��'T�._�6�qӺE���O`AB����KY��\ R�톧Hr�����~�j D��1o���H�}���O�lP�'a�:DR�4P�! �	� /?����	��?�&�������?�'�?����������˂��,���K�r���A������?��ih2l[�y��'�L�ڛV�ǬW���!�Ϛ'�R����� H%x6M�=~/:l�����E4O>p�bן�u�4+���'q��1G_�b+̭jZ�����n�d���q�pa�!��?q��?���=V�i*�.�f�_�p!�b����Y%i�kz��6O��D�O>���T��I��M�;6�.@��pf2�2�̝�$�R�`'�i�F6M���d�=ܐ��˟�(�ū�q���̎3w��z2D�;��!�7�X=('��$�<�����O�%��#@`yL�O�;�ʧP>H��̸i�еbL�1^^���Q�Q��d�O����OP˓K>���w
T�<i��?��b/�p�zE�F�$��U8��ԓ�?a�Y@~-�>a��io�6MH#0'�$�� 朣u䏡N��ԡ�Dߴfz���فVx�`H�	����m���_>�6(�O��p�����qϘbBt|@&��N�h[���?�~ǲ\�΂����?���?AF�Ě�lM �Q�O7�e��`��?	��4�H��'�7m�O ��3���]/��u��	g�\j�Ă@G�����<���c�4NLNY�B���u�"�|��dӍy�L zZw^0u��L��	����aA)\~D�4Jm2��'����̉��-ځ��O����Op��3T���e�F�<�(퉗�P-h˪hCvo�<A����_�<�̓�?������`~�"0=������f�^1Bu�*I��U,���uӸp���Ox�P�P����+rb��C�R�r� ���C$�� �@/>����0O08s�e�j��S�%���8B��Ȑ@	�,�6@r٪d��1bhQ!F�]0�ZM�V���\:0M�� lH�š�+�/\�¹k��+Vv��`ţҌ��*TH5zv��	 nŦz�� �׎Ԋc�Π����u����c@��H�j�1y�j�vH�?[Cޘ��O
5D*�PR��Jü��0%�� �V8ȕ�Y���|*O,����鋞feD��M̢(�L�q��A� |4��� �D~� ���I�@�h�@E��6 �e��
�7+�:y����M�%,�9�`n7
���%�n��@Dl�:|�2t@򪌘%�p7�m^�$�O=��O�T�'P��;��$8�vD
p�D	=��9E���(L�I̟��I�@�'�$I�~���؊Ay`�ӀG*��&,	�
��a#�i����4�~��(�?y��U�^�{"#��u�$Ģv���$(�����Mc��?Y*OXݢ��z���'��O������Y������C��<�&�W7�~2,]��?������ۋ
o޽�7dN$��:�F�95���Q`yӄ�v0��i=b�'���O���!���'��z*$)c��M�# 陥K��?���a|�])�����' ��$�T ��H-H�b��Wx|n�l5����4�?����?��'Z��/l�&牞$����@F�:Z�6 pՍ�Wnf-��4#Hf�����&��|���H�[ã�%~\ݡT�֬ :h��iF��'��i?A%��%u����?1�nݦ5� ګT�M��F������
8�ɯF���&���I矈�Ƀh�� ���B:P� Q�1��5�ش�?��XN=�	�f���������i�����2��RƂMk��+[�`�$�L�����%������L��Hy��+9$��!�[�,R&��~q�`-�>� �B�<��z5̅��?��IПx�!-.�0�2�\;r�X�n�K��&�p�I̟���iy¦� �	ۉ0�	��	�T����}w�FFǐxu��'��-������?I��6�?i7`��r%*��6F?j`��3%N�g_�������ڟ8�'YTs�,�~R�r%2h���w���!V���<'�8�ĵi��쟬�~B���?���c�X��{�
��	�Ǝ��$v�@������M����?y(O�E�1��O���'Q��O�z��),+�`��J�N�4@cJ��~葫�?�[T�،"Cxޡ uL�f!D!�Φ[2�Pzwvӌ�/���d�i�`�'�?��'=e��||�-4V\ҀKB� �y��H�C�~˓8������?��yʟ��ȼ ��}s�`S(�L�끮�M���8͛��'���'��DϹ<1�~>�/[\��PH@�'3�I �蜯mD�LoC5.��	���'���<�������@��&� P��OݫKZ�X�i���'��T-;���$�F�蟠{�Kv�4�B�B_`�[����k�����ivR�|b��~��?����?�BG�� :�Ï%	OH���N"5���'lN�����<12�j>��I�4��^ixWd�v�uZ��޻-��@���xr�'p�'��s�X�I�`d�a�M��HҐ8�⋗b��tb�'QyB͍2x]�=O�A��������ʙ�Ȍ�"b���*��&��MÄ��f��?�-O�����~�z��7�l��a��dX6�(j<�m�0������<	������Ofʧz��EnڸZ����sY�$qc�U`����?i���?!,O~\��*�W�Ӗr�*��Ů�07w8H����k�rԡݴ�?Ƨ�U?i��]y�O~2����L"3�e��̱%LJ�c�\�����'��Iß��$g�Y��'���5FH�2z�Ό�J�1-tνI��3u�D�I!(#���m����`FxZww��5o+��p�p"X�F���4���[v�%l�$����O:���ByrE 1�:E���L�vp�G��1��/O
P@�a�O���?�)nڼB�>����hy�8�Rd��k��6�K�d6��$�O��D�O��I�<)"��|*�!�B2�@���"Dd~���Ԕ|NR
ʁNG"�Ex����'�J%�dB��j���w"=2�0=�`�b�>�d�OL�Dx�|T�'B^��'�?�a)X㦑�D�  1��0F�J�
�d#���|�$"�D�O*�OR������0�!�K�3zEra�P-�c��'=�q�P_�tåAp>�͓m�������;h��ec�"յs�!s�^}����?����?a.O��8�V��@`��^�-�.�Z��Y6�(�'~,5����?����3���O�S�)d�٠bY�9B��k�`��7�O��?����O��`p��?-�Qg�6T�F��"J�i���0w�t���+�"�O��ɪ5���O�"^>��B�x�����ɩD�����jK������_�,�	��\yr/�"LT��}*T�%T� �2!L�m��-	E������$-ɂ�ɨD���|z��?�Oj ڡ�۵:J�e)��O;�q�4�?�,O��$Æl�˧�?�����s�9��C�N�D��llj��C�O���2�'z�v�͈W8�ӺBF�b|�� uҀH�4���m�'T�X�(bӪ�O	��Od$ʓ�@�A��IQd��s"mI5u��D�J�^y"��H�����9O�s�� �ٱ�?ځp �w��I�ճi�H0Sp�'ZB�'���O剻Et6瓎mK�y�,��0g�L`�	ߤz��)�-���i7�Ş�?�%^�+B�Y�sEɚ�T2���u�f�'zb�'��{!��>�I��<q��  em����p0�͓�(��iP��ө7�06M�O�˓-t��S���'2��'��D:Em�M�P�aR
�JZ�+c�cӪ�dQ%@h�L�'�\e��'��D�y���5&`�0pd	J')��h�!n������~�d�O���O6���O���zT��LR����K�s�Aː�U��	���	П��1Ku�������I�(ʴ�q"�^�x��5C?
4��D�u���'���'7�V����吐����Ǭ�&H���U�(�h����M�����<A��$2��������?�&���<�UCʃ���&��L?tP{@��������П��'ՠY���~��x�C��]�q�ĸ��C��!xJ,)�iioK��y"D�'4D��'5����O���<@�|�բڱ��X``A���6��Ov�$�<��"�0TJ�S�\�I�?AI����_�r��.oDZ$�'�>l���	�d����	ҟ˓�d�&��c�w�n-
��_�G%���& ��^�`�4���Sb��lZʟ�	ҟ�����DQ�B�$m臅#ϒ}�qGP0hU(e1�e�O���Ù ���2�D��ʉOOM�b�N#��1�e�V����4v������i[��';��O��)AP�ϓ5V����Ȍ>0f��!jUn����i�:(��'2�]��i5�?�S��,i�#
  �|xR����!0L
��M���?y����]��[�xj�r�h�ɑ.7͏�"2�ZԩJ�7/0U1f��ݴ��� $�S�d�'��' D���)��^ypVႺ6� @�u�>�D^�t��Q�'�y��'���*�y���5&�|��bp�΃7�v�� X���D@�E��O��D�OZ�$�OZ�@���.�Wd�3/�ْ5�۬X�X�O��'?O��$�u
��n�d�O$q�֨FF���x�"]+5d�1*RjM��������Iџ ��]y�䙵g�<�SN:��S���R�*��ԥQ�VR7-���$�O��+�8O`�i�O �$�]i�	;�*p��MγP�䰲�0~�6��O����O:�ģ<I5�o��W?U�I�
Ѥ��B͉`9 ���k�C001�4�?���<)��Q1�?Y�cO����4mI�E�O��|��|�e&6(
|m����I_y��>$맺?A���:I����r�Dڵ-, ��-M�X߬L͓G�����?�%'�<i���DV���c/��?�>���
�:������a�'D��+a�x��d�O<�D����'���S�ʭo7�(��b^$�}j㙏e�b�'��$��E�3T�'0�0(a�&x�
�G2kXڴ�4 �Bt�4�i��'lR�Od@�do1�%��YBEZx�dH�2��	����i���;�O"�$;h��|"�7;fHX�*�N�ECF�C��� 2���'���'�8ܳŉ�>�d�<)��G��toZE`����.����O�?�c����b$���`��ϟ����Ɨ%�4�v-#t������M��ED.}��^���a���əK]��I�?�+Q+D�j5��7x�Ps�Ǹ^x�7-�O\ �50O���?I���?�+O E�.�xP�H�F0hԩ�'-ǳd��T�'�&=�'X�'���y��O���'�R��������%Uzz�4p�ꛑ��D�O��$�O��$�<y4m�>#���(K6���Y�
���v�P�I�����yB�'Ú��'��4�'u�	�y��vcDi �)	1((�m����6M�OR�$�O����<��W�l���طI8�;1.�$$���G+E�qG�6�O�M	�7Oj�җ��OR��֐S<�$6}�)��s��D���]�d�Ո��S��M[���?A.O�REy�S̟@���s���G

7�����( '%�"���
����ծ�O:��) �%�$˼kڄX?��J��xG8�p6n��Mc/O���[�����J����L8�'C�lH��)v	�F�]b+:��5�;�?���~�<ɶL�B�IV�@�`�g�z5Xց-y�(7m��B��nZ�p�I�������"�yR.Z�+�x���/Sp��E`�N7m�1���.�<\(1���<k���O+1�Ay7%_ wL8to�۟��	�$�d-9��ܧi���'�t|��4�H5`��4j���h���?_��EoZh�q�:�)����?���RҜr2�D�88��6�6Bq
��S�iJ���,a*`�f�<�	��po4��sRM�B��,X�S��Y�H��':��t�'��	���IC�jp���԰;��9s��a�����U6�R�'o��Ο����O6$�&i�7.}�qq����
�<�L���$�<i���?Q���d���L�';3@�EM�=��]X��̢kZ�1��	.P�$�O���4OB���O� u^��d	 ��}����	�(�A0k�QJT��'���'��Z�Dkc�ħh�H���D�A�X< ǅP �puQP�i>"� �~R�ڨ�?���T|�����	�[d� a K����{�"6�O���<�l@.F`�O-��Ot�hA%h	�x��9 �d]&dm0����~�Ǿ�?a��S������-��%l5P��t"� %ظ��r	[ac��]�`r��	�z��h�~���BpY�dX�U�r�Е� ˣIdD��eJ�TfR�$�OXHb� �O��O�<Ct��䅅i�����l_�	Yt�1�?�e	>�M����?���0Y�����O�Hs�#X� ��P�D�8tf�b�FȦ�ba�u��'� �u�1��̟��5m��X�:T��(֝V6��v���M#��?�����1�P��`6��O��䒫���/\�t�*�*�IJApUK �]��M�O>Q6�-0�O!��'Y/=� &�{kωN|TiR 	\�<s�Ux�inB�X��&˓y�X�S�<���'nZ�Lfލ�Ƅ\���UnK�25�O����Oh��O����O��"�Ԩ���Ç?-���ҴIZ9Im\��	G6N�}���?�Iz�7��2Q�eZ�i��ٮ��)֦��	��	՟ ��� �'*@�X�~�΄`7��(GP!g��=�Ȑ��i��4��'R!­�~�'�?��jB���Q6ɂ�#�Y��a˗p� �T�>A��?����DߴK�a%>A�P�R���(�.��&�ш�F�8�M���ۚ�(z���	�<����1c� ��G�L26��#
�X�L7��O,�d�<�٬HT&�r���XAH@���"i��\�%af�'��K�ćR�"3O�g�'oM򵨉���TɅ�DTH�4��dɼ#��lZ3��I�O�	�NyҥG9
�؉�"\�0b6q� BF�`p-���?�iBW�'bX2I<!�� b��`O��Gn�U`ƈ[ڦ=�$��MK���?����BDV�����O0`�`���']p ���;YҙaF�٦�`	!�g���<1��F�^�H�n9~S�qC��23o�����i+��'�oʂHF�I?.��S�XY��d��5�T�ܖB�(�[��J,F��STk�|�'u������O��DS�E3�|Q��S.0c��ӌȤ-�Tn�ӟ�����D1�i�O�@�`�h���ihha8�.�!�U���SFB x`L<�H>����?���?��m��0EeL�&�m�w�i	�¥��7)^��	ȟ�K"	��L�	�o�f����Db�PQ"B]U
���F��]wl�UM�¦UPT�>?���?����?���ܑB�O΂5��
Gv�m���%�WcӒQ���Ot��/��O\�3O���B�M��iT�;�(�! ��:�Pu(smL}��'7�'*�	uH�!ꭟ@�DTwz�}�u��5�@GF���o�ޟZ�V�<� �1?1�'ܸ'P�-���*�D��C Y�P��USڴ�?��?���G���J��?����?���l08'�5�������78��1B��O?����͓�u����O��U*'���!��w�`h!�`����'"��(��'J���?q�'N"�cむ�8LbQa��~#�dywJ��@/�4O�P����)�O�O�,�h���
P�<$�g(Z������4�L7�id"�'q�O+@�b�rq�'�dqQ Y�⅙�g��<� /W&{l�ւ�2�ў'���	F+Z�A�@&7.F�0aBNB �)�4�?���?Q�m]��?�L���Χ�?I���Ʀ����9k����6���(�r�C����O�'>��	����I>R|���ӱ"nfL�VJ�"�Z���4�?i��_��?���1@�T�'�?���
Y?��\�i��=W<P�@��ٵ��M�K<�v�L~B�'���'�削|���Y��q���tJ�=r�i�*�'��$@6g���'���eU>�MܴsrL�JC�\�h�x���#�o�h̓�?Y��?���?�T��5���mJ&\Š��%�L;� �1�$ˁ�M��K���?���:���?��I�<�>1%X7� =�V\�w�L\�Z2nH!��I��?E��[�c�<$�� �[H���&kP.�y�g��C xp �M�tq ��:�~R���!DpB'���#��鸳oP�	(H��E z����o��-�n�Zpƈl]8�q��@�%�6D�g��s�a^Ql��!�L�F�����P%���M��������'+h�3�C$h�Α%"}4`�"F��4�dȷ�7W�����6��P��Ι)H�л�NG��?���?Y�he԰0�`:{ߦ��Q�D�M>����I�#�ά��@E�O�d%=G�YN?�DO>�j���;#��ɢf�!�����[�'j�!2��Z��)��tY���X"�� ZD�IهAFfIЁ�I��䧹�{��9�@�	XlQ�U��; (jM�ȓT����Տ!fH��b��ʷ .&$����'������O���5|Y�i�G��e`��r���@�:�D�O� �W�F�-����OF�D�O���%�û~`h�d )��㓇�$pp�躳@�u���ɭ	��s��+C��1�؟ў� V��?�8��� ?W�ި{�B��?���?crLB���#7E�3�~���Z��A0PY%L�/G4��<̌����F{�[�4�G���$����eR��d?�On]ΓQ��$[��R�1'Px %�P�)���R$�A��2�'{��uāҁ
��F�KA��i�&�"�OY�N=�(�I��t���<R���6S#"�I�|�P��A\>��c9-�*9�bd�xL�kю�"$���(��<�#�����⍖&Y(}X�_F�@�3p��.#��iQ�_��<	@̟4�	-�H`9⡈3�
�%'���|�E{���-��h0,�.� �Qj[)��#?)B�������J��3�DزfgG�-�J�Ʌ5q��ky"jA�<�z�'�b]>����[��5�Ӌ�%��jTv}�U�¡Wǟ��ɊY�����Kώh�\�����?��&Ӵ$�	�zw�@i�JJ�6��@6M1�L����růIW&�`Pl�<��'q�
	W�
/Q�vT
aE�X�)Dy2��?����O��C`g[P�J,
����8�'u!�Ԣ_�@X8��s0�y	�gĆ����_����~��	�e6԰	��G�T����f��xH��I�6���B�E�̟���D��aϢG3R�'<��ɒ������L�lh��h�!~�E!b�ȓ �`�RO��I$�S�? @�X�B6���Z��Xۂ���R��"<E��{R�\�o���Y3Ej�/Bc�m�W%���?��y���'J���kC8C��9Ӥ�6K����'�
A"6��U��Dq��s4JK<��8O������	* \\���_='{��t��#�C��"G�.�
�)�3q.Э�)F'$gbC�">6�9���:�A�qj�+�nB��C��S��O�#�X��q��p,lB�ɮ}�H��
�v��(q���:kjB�IQs0�0�b�pؚ߮f�I�_;"C�I�M:>���WbZ�X���	���B��8-�P�ĄO�:ǒ�d�ўiw�B�ɋ>C��W�T�%�nl�BĐ9f:C�I3s��l`� �<�JȘ3�
�R� C�I�;���
�u�Ҙِ��MQ.C�I�+ư�đ�d�� @!���C�9'�d�p�=p��SPGԝN��B�	�!�%�Q8�pkp��2*��C��<c
�ɕ�!�*�X�Ϟ)��C�	�	��}�A,�'0h� �T��B�	�:�28�Cƅa�Hb�� �vB�	�=��yC���V����ŜzZB�	;H�����H���pB�6��AvG��-�0x�nQLנB���ycd%�(a�,� �k��f��B�l�4�ĩDc��@/I�8��C�	)W��
.��n)B�i��� hVC�	�DI>q�PE �BU�]{¨�C�	?zX�CC���4h"A
>2JC�	� A��lM�<��d�c�>n��B�	;���{�CC��x�׉��w�~B�	x�)��d�J���H0��%) C��r/�����K�@��ǣ[j�B�I�^��0!��Lc5a�+H.�B�IA{����!�����C���<"�B��;�j�#!��'o�,� �HxC�I6X�꼹s��#�z��aS7^�B�I�\���q�N�Z�`Qā�p�B��/wrxȚb�>=V\����P7��C�I��=PS�L�]f�Z��O�όB�	�M�.�ѧo�$L^�BUK�xB�?^��qQ�۵W}^ͪe�;G4&C��/H d�Q�5�ꄩ���� C�I�����.P�� $N��B�I�b|&|�dƐ<tή�j���,�B�9u3L!�"�AX��聈|nnB��"i�թ�@�?$"D�a$@�t�\B�	�$DЈDG^,d����3��s�HB�	'5!s��#7K��y$"
	sB䉐J�pEH����E�4Br�HB䉫g������/��ih#.L�	pB�IS=��HV���9�2/`�B�	7��4)�h�GWd,�����G,C�ɣ+�Vx)�Hϭ� ���o�*�B�I#PT�w-�:W���w��(��B䉙4ov�!�A�_����p�B䉒���(�L�@̭Y��Y�Z�B�	2a�ae�^�ݘٱ���y*TC�I�1�ʔf�>o!<=��ʖ!A�:C�I�u�|
ËЧ9Ӵ2��E�A~��m���M��g��G�OQ>�iuΛ*��qKS��0��#�0<O���KRm�	�=��p�䄖�kOR��TI*�OB�����<YG	��� 1�ϬOr��Jg�W���]�� ���De'��'k~�H��`Y�=����d�[H<� |�W�¦?��-'* "��� �	"&�=Y �Om>L���Pܓ21:�C�������K�N~���	�'ԁc��D/j=Pɻv��;-A�QR�	�B�\���4}߾�:'%)�)ʧ����QkK>B������,���I�)�Y8�?�D�>A$2�b���.vI��+�;$8�'fi�u+�yX����ސ](4�E͙a�Mِ�&}��1%�xڊyJ|�q"R.�˖D݊��X�D��J��(��:$�$`W��e��ʆIL�N7��&MB@̓J?���M㟈lv@ٯ�'LN�AH\��`�䧘+HxN5��OP���_�*5�h8}>8�KW7$�`���i�-���.�)�'^���s��}�0�2,Q�J�d�ȓE������[$}ժJ�G��Om�̅�T��-��pW��y�F��J�\|�ȓ.�HP�u�,{���`������%��	t��{��L>����$_�(H�J�50Q���[(<FbS+V�D�1 -\�)�z�ڶ�Æi���"�M�����d=.��/֩�
� "V��]���Z��p<iЀ�``H����7?I���i��8��e��GA^��N�v�'CJ����S�`�����f���Dʪ3�L�'��}�1/��Qo2���2|��
�욌;���HA N5I �I:c�t��?E��fV!2�ƌ� �Z9�~��J��7av5bK���U�gq��'
�(Т�U���R�V�fQ�)BJ ��,.pҧ�� )<�@×�b`Zb�$d*=�!���8$\y	דA|�xӪu��@ߡaw�I���l��< VT��1�MT���D�	4���_��X�`k�6:�f]�A�&9Q��.�g��U1Hz:擀W��X�ā�;�e+�F�L�bB�Iz��q�À'��!1��/�N��(I�O^��k9�%�����r�J�р�[&`�ʔ�ȓ��Ë����4�c�+7ڜ��I<5�h(�?E��/Υ��4�h^�� êނ%�!���4J�b�ʖ"ӻ'�䀚͛u�!�d֜Cf������y�99Ӈ��:�!�W';��Yq�B߉Z���Kt�C>�!��3,Ds3���P�N�!�$[12��H��8D�p�J���W�����"^�=*����<�hҠW�Q��}R�V�U��d�T�`i�1�C�	���$-	\�!���*�ve+�L#`��b��=�ў,¦��q�OzB��H2i�Jd�S��9[����'��e����'r���r�֜27�))��O�\b����~x��3�
�8冀��BJ�p�B�ɋ3����b�#O�zlR�"e��˓�,9�	�+��}�#Ǘ2y֍P���bĞ����f̎1�
C6��s+ٖ^�0p�I:6=�؅ȓW���tK�6$|軣F0~�MD|rJ�<���R���e��y��C�6��$yb"O�(��*��=�>|2`h�9d�z��"O���0kԐ}���T�<8����e"O�9��Ř-t�90g���oa�DQ�"O�T�@A�4EEm�)αw%��q"O&X��/��v(���� 6r��	�"O\|�AJO�z�m[�Dp��5�	<(FƄ��Odh2��)$�k�MȜv݆��
O4���C�z`����$�k
��a�'��,��No�	�	�<�G}"�+{L�Q�2�.^S��`����O�0+C�ۄ'8xL���~ʢ���4�V2 W�4#���䦡!��p���ѓ�W�yd2�!3�"y"J�"�Ʊ<� ��04�*�{~Zw䖁�G�O�S=V'�tgŊO.� R�X��B�	
Mn�$R�%!H�q�ݿCC����^�@���i���{���Ĭo��4�hs�ȏ?Y8����@���=h��'��e�M�Z'���W-�3m��Cr!�&q�����x�8aԦXd��<c/����S%zݵ�>a'*qW
��w�}��$W1
WF@E|�FD*pb� e�Лx1��(F��(�yr��`�8 �F�&oB^Q���GN1	҇�(Ԏh���W�����M�7En��c����6�B�Os�xQ��YF.�L�ub�D}4���E?��50��� ��I����� �Dy�"O���Jѹ�|a���w ��IS��?9��	���wܓޤ�X�5���Pf�+�w��&,D
aN�rT��N�P��Q�ʰ-�DI
���m�!�򡋣N�M�+O�=(�ڧn92��B@`ahˡ6��c�(XV�<�)��'��8$�=ړ6��T:F	_�7ʼ-k�Є���Ts �Zp.�	���PP�I�,�2)B1P�EgR��ub*A-�5���+bYl��k�tZ����l��N}6�DІ*<6HC�YK���o�"��L8�$����0k�Q�+��yK�AR�z3ꙇ�!ޞY���L9tmb,���(�n�����#<��iě6h��ZfG�%���ڝw�]2�"��$�x�um��7ט�1�/D�9����+%�Q�� �tQ����4Kc��c�bMY1JMH�YXM�0nV��pӐ��2j�Ɛ�7攷Y�b�a�
X�">���:Vrֽ��#E�%���"G	[�%T����3%�4��=/>���K��x"�8����d�wz�aڰ��y2��Z�6�:#��I� أ"
�Lk�����I�9e2 ����0h���4���V�!�^�~����",^��M�� � :����3�^nB���˦;�-��?�+B�v�I�O�|�z�I�8��lsg*lT��	���\:e�G�	ǜtq�-
�0��ХB9G|j����X5^��	W�H�L�*���ɡ%o�z�àN��$0s!T6ݜ#>y4�� V��AXT�؞@�.�Ʈ����-�4�/oF���ʀ�y�$jCΐ	��B�?u��@�Z#`$R��)��*|��	�JY�B�"���H�Ư�5R�A�J �q���f&Q=sX�PR��R�e���B�"O\��ɋ�?ֺP�eǹz�dc��D����g��"�f���)@4B�S����xן>)�k�%y�|bt�Ր+>�L�b��ؙ�P�X�.���EQ<60(���	ˆqᨴ���S�!�R�h�m�Z�>��xZ�3��{�G�,c��y/έۈO�p��f\�g����섲cO�Ļq��X��3����d�)�!�u��l�ۣ�0�LbAc@�=<�1��-�%K��Vr�d�C#1�x�0d[$� L`EkP�}��0����*XoG:�1	J c���%����yRǮL�@!BVj�x$-��O��<}`�Ȱ$-6���HӠO󄹈˟Zmb��!��T�+&�ܚ��].X� ��4(�~�a~
B�`��|��[��d��!ug���%^8G�D��0��>	
Ps���9�℅�I=D��b��C�Tn���ʯ��">���V��XH*��q0@P�1+��: `��>#�ٰ7�shT]��>��x���:b��W��B�]�Ѿ��'W��q�g߫;��M�ANOU��N &�C/�4��t��.	���܅�PwB]@� C�DQ�9�v��0V�<qq/�%d�2uKM�#�y��W���dU�y XC��%4��9�K �t+!�&Y�Yz�)�c�r���$ J!Xi�1鋅�Y2� ��k����$�0u��B��   �
Œ>��z�(@�2�@��� Bx�#��64���s)̂X�H��ʇj�<Y�O��K�!Z�E؉6?�4� M�@ܓ_�|��M�>��]�� !�'u�da���B���D�\��n�f�<A��de��F9x����i�!򤈩U{�Z�ɟ�����F
�t�!�D�i��ěFoۓP�x�Fj�
�!�$�:r��X�T�DC�A�u	��i�!��^�,����\�~/����%!���-w[��QtS?C����̙�I�!�$@�Ph���R��"J��!�d���ntQ%�
t��Qn���j͆�S��p5/�(R]*dc�j?� �ȓA~�� �3c�z���S)��d�ȓwg��*%N�;B�<	`� X�Av���m�6��4�0h�L�CF�~�F|�ȓiG<�)Go( 	�����U��Ąȓ	���!�?AN�R�T[Yj��ȓ4�>1�e}Ħ_#(R��iQ.���Pyb"�%rV����J�V�|�%�q�<!�	�C���'�	z6�(K�x�<!k�2h`���W;F(���(�t�<1֠�!P4J��f�K�)4��x��Rf�<�6���gUmpQ(u,_�<��`�pk�i�
���  �]�<� ��i�HJ	�r�;ԯޫ\r��P�"O���D�S�+Ր�0.�)z�ڀ!V"O�l;��5(�b��}��(v"O��Z��ֳ*d�0[��=Tؠ9� "Oؘp��AO�|3�n���q��"O�:V	
�clZtx����쐖"OBə@�=3�~yQ�j�'��H3"O�|�W�� &@Ԋ#I�
Qc"O��1�N�X ȑ�<�L���"O�P�0�,yLB�K�1Xb���"Ot�[�fؖz�����ޯB�� r"O� c�cI�x���&3�����"Od5��(R#V��٤��#F�� ��"Od1�4b��H����MP���IE"O\E�cĘk��1����m�E�"O��3ѱ>�@$xO��43�"O�;�b�-2��3��XBd�7"OV�P&�O�I��7"��].PQ6�0D���h�|Dد���[�� �y�CB+{#�-�@�V/+~܍Ё���yR���(��'M�*Cnh��FP��y2g� X�`O�6lf\�w�U��y�$�<1Ȓ ���#B�(���A�$�ykϥ7���cS�Y��*䳇�;�y��B�¡��!s�p�giݰ�y"�][���!j��$j��V�)�y�8y��R���sOF�R�Ƙ��y�ID�d؃�	� @'H��M	��y2!�N�D�AR�m��� �P��yr���CK�r�.\�G�ѿ�y��5�~�+4(V�_�I0t���y"&$M�� 2�N��P�6KV��y"�*�=�Z�J����Ѱ�ybFΫI���r��.5�^y�v���y��X�w?���e��*�u+�I ��y2�ߪ?In��DV�&4 I�����yr-�$��9x��
������N��yB�V�OXUҷ�D49�܊�AN��y�"�sLK��Z���ue���y�F�<"%�Ţ͑OaBYp�"$�y�F��x%��r7C2R�V�5M�3�y��&F�=�$.�J�B���"�y��<WԼQ�nQu<ur$�Z��y����jتvO�4OCj,��JI'�y2K�츢1þK���S"���y2&_"v�^1�5���J�}
����y"�%HȔ��@!p��(��g�)�y���`7����,�u�hy�g���y�k͢t.�т%��8}n��w+���y�/W�[k�1c���
yZ@�W�ݵ�y���FŌ�bM�l����v@��yN>z i�˱aU$ղ��^.,�=E��IE��(��
%�&L���4(�*���d|��X���"l���&�r���ȓ"���Q�E^�$��I�9�0��E�l�j�#@�mY�i�6.B
�����|N9�HۉS��m�fgȊ\��X��;�,�:d�W4SUxxiG�F��%�ȓW!P([U96ш�
��ڞń���\��ʘ�$���$ʿǦȇȓU^LyH㎰��M�����qRf=��w�0��.��u�4*���Bm�ȓkQݨ�	Q�0"$����5wZz\�ȓf�P�%�,i�2A0Vl2{0�M��S�? |�h�n�&`0�"��$��Tq"O���bR8jS�!�G��EJ)ض"O
q��i�6��ȸ������"O��°��[ >�@ECX+g�J-�"O����E�P�U�É�V��lz�"OP���$]b�a�'��{�"OV�G��)���0��j
����"O8Aǌ,v�6�����WW��w"OГA�U��K��
j<���"O�y�� 0�|�lJ ,�)�$"O`�Ы�yI�A!%��o�μ`"O�x 7I�+9"02��ZP�����"Ou��E\!($ȉ���Y�)
p"O�����K�$���d�u~R�("O�i$G�RB�uq�柽�R�H7"Ox��Kځ�f[r����0"O*� +Gvo�A����K�f�X""OTM� O�
����B� |��E"OL�y$�� ��us� �]����"O�3ǎُ-)�������h""O�@����A� %�q��M4�!g"O�5+@�֠b=� rA"$-Z5��"O��1S��E�eO�[+��I�"O���W��$���;R6����"OD�de�S��4@S�G�!�����"O$��$�
,��K�45�J8"O�XSbĮ!�Fay&��/� �C"O� #�dV�Bm}P���;|�p�(�"Ob�PA���$��Y�*����%"O@���hǣvS��D)�O�>({""O.��������t��'j)J�����'�ў��V�ţPh����L�0C����4"O��3O��Y���q׫�0x����"O�"g-��x*�i�Ikh|P"O�H@�$~F���/�/��u��"OB݀�DB(
l�@g�>����"Oz� �; w�a��̞+� =;`"O���vC�*p��]YY Z��]ғ"O�r�kMt�p\�"H�:}4E�"O
A#B[P��T�f�k E"O�$�<�`$��e���H6"O��)AØ�m���6��_�N�47Ot�=E�$�T�8�6�����7#�Hat��4�y�AT)H(4a�B`�&Ͷ�k�H�?�y�ā�]ʘ����S݆������0�S�O^Ġ�K�/G�`�E��{����'�P�Z ���A�[�h�J�'ΰɘ�KWvm��DE��|��'Z\�6bR
�v�*�#��N��`�'�H�QC�� ��	���~P�MP�'[*��A�Z$�WJ��}��}��'�X4)񊑶:@hgB+nS�ݣ	�'�ѫ1�	�T �
�kRF���'i���f�7L���k"	�(j)�'o򷄠K�r�EJ���M|=3
�'��=�b�/i4)+u�ΑA�i�
�'h�e�.�]#u�J8'ytR
�'༸�KV�
6�L���Ζ����	�'\B<�!
��E�Q��:Q1��'�l	�S�uF�)0#\
%y�
�'� Db���P�R5�w��
W2,8	�'Ƃ�+�WM�V���%�	�'{� �Kɂ,+&�Qg�).�@�	�'���3��}".�)D\
F<5(	��� �x1wm�#8Nx���Y�b��"O�	C���F`8���.I��7"O�TS��z�lL��o���H#W"O�0��ܾ'���Y"�ϔC�49*S"O�¢�jP��ۃ�OQ�h���"Oƥb�OwԒ��t�$�:���"O��C���U>^����r�x!�"Oؙ��]4$���#j�9�� If"O�q:�#����1�Lk��H"O|�b�,��<]`m��r�{T"O@P� !��x� E�g3X5kw"O8҇�"vƶ����@����"O������$f@P��	I!��A�"O�(HO�� �pd�ǁ1UV�E"O�Ґ�ò)���x�g��w�H�"OV�!��T-c��ᰈA�U�`���"O�5a O�4d�t�]�e�ҡi�"O�����Ev:����@(W&8#w"Ot���[���ՆU&.�Y��"OTX!��B�T��1�ȴ'�HQj%�>�����~��G��I�e��Fw!��ͰQ���p�^g[���f�>wi!�d��; �tE*lzTՙ���^�!�$�&౸g'X�r�x�#B�8'�!��P��T��
�gS>M�!�P!�D�(�d�e�&)4&qj�B V	!����3�4�Y�-$���"O�`1����mK"ǋ 
���"O�"t��"i�m�!�L N
W"O
D�-W,:ȶ� �,�"	2�"O��cZ'S�XQ�Fō�!��%"O�4r����Fr�T����,�&ѩ�"O�eXEO�Fz�)�� '�Z%X�"O>��BQ�l M0�LY.5�U��"O��� C�eJ�]
�r@p�"OR=CE�X4�ذSPʓ*@�rE�U"Ob}�e`�H��Ta��Na2m�"O�A9�h�"���P'�4k����"O^�{���8X�F@(#[?����"Ov4��V�R�� �e��zp��"O�q��̌t`���M�i	*@`"O� ��kӕ�8�͇7�>IH"O�l����*Y��q�,��G�L��U"O�]H���^�����c���A"O�Lڒ�E/ZaWK�%l�B��"O�Tq�k4>�ڡJ��H�${���"Oj� ӊZ2�����+Abe�|�0"OB�*2J���X��+̿dFm�B"O��qE��A8Bl�UIK-sx8��"O")��k��/��0s%�g�l�sP"O�����B B|�$_�O��1@�"O��i���X���D K4�  "O��ɀ�\�NJ�ys�!�7
��"O�����7=�@�p���H��)�'r��۲��-�&Բ�.��
v4�h�'�>���b��.�T��U�n��'?���� X��,�j�:�d�
�'����B�r(!�o��ߎE�
�'�pᑧ���
u�U�^T��IZ
�'�`���cuR�X���JNhY��'@*a� �՜���%C�\�U�	�'\��+E��U��P��=W,Z�'lƬ[�Hۜ)��(��8m��0��'8��Tc�:Q�L(CcIhK4� ��� he�`F>L1B�+C��(�"O�l����(��Pzq��,*D�"O ��Q5�4m{��,,�J�"O�a����� U~a`�Jq��:�"O����BR>g <Y@�k��b@���'�l$y�'��Rv���i �C�0���'V�qPؙM.ƽ�1\7m�٫�',�(�e�iY���P
��fޜ$��'�� �U�E��e�K��(9�'N�\�A+���H�`��q�:MI�'�UX�N.:+h+����c���2�'�}Xqm>x�@,Y���W�<C��/�D����SJd<���t��C�ɓ(p�D{���g.]��ׄ'�C�ɧM�ܔ�(ZY�<���*J"�VC��.�8=I�
F,�H���'a^�C�	���0����}8�@"��"�C��)KA��a������ъH9%a�C�I<o+�� #%\*!���q^TC�	�+J�&eR7j��s&'N#�B�(Y�2p`�,�]���
9��B�	:O0f�+�'ťH�؄ �	,C�VC�	.!�Lq��Y�4a��kU�Y2_1.C�	<e6x9&�ԯ|{�PPp��
��B��$l� �����l��pۦ�s��B�	.m������o��dk�2TC�ɎV���S�+�#x�X�,�I
C䉇\t�1#Κ�{�޸!�+N�4B�I%`k@��엊%���+�m��.�hC�	Y��)4�B�ڮ�#�}hLC䉆}�lZ��]�
)�LB7��9�C�I(=�mӓ�U�D��(����W�"B�I9X�۔�ʭ`�jڲ��6R�RC�I:1�4q�g/�=�Z� �"�C��>w��A�k�(7T4�r��S�V��C�LQ��[�G�*_�\�qr�P�2R�C�ɠQ9�� �g� !$6}�Uh[�6�BC�I�+B\y�
�>B��Ą?'��B�ɟs
�\�Pʁ	 ��$M��B�	-9���1�Ēr`��.�5>ʤB� Rʤ�'"��GD�K1b_�^lB�!r�n	�#�ɫJ��I#O/j�8B�	�B��Y��P���X���*v�\C�	�|m�}��A��F9b�(Lv^B䉆|�0X� �5�"��@�
'�:B�	�h���D�d�`�bH�2t B�IDC@m��*�{�l�r���qhVC�	ZkX-(�q����ۍ%aVC�*\�`�2�B�*�>#����|*C�ɬ
��zt-�-�ْ��5d`C�&2nX<㱈��CaҘ2��KT`�C���6T�c�րnP�<�� ��̞C��-"��1J!4��dz�"js�B�I�EL�1���eɮ}�����B��?;�z�@d״-�891!N�
�nB�I�p�d8��=��ձ� �2�4B�I�2z``�Ήl<�T�w�S�N9PB��.lXlc�kW�,W����N�|XB䉷)b���	�1�p,JP�_|	LB�?��d�!�E�v��� cO�B�	�	Wp�ڹ=%�
H	&C��82�G��%&�Ҧ�C�ɷ"�[��Ǭ��2D�nZ�B�IiQ���[��0L�k҃	�xC�)� ,u��j�$� C��8Y��Hbg"O��+�@P���	���)���G"O���ᅼΒ�ʑ�R������"O0\l�n&$�僙O�A�"O ����_nҾ4����tM�3e"O"�a�aB�oSFy �oX�9g"O �i gӻ@ 2x�NQ�~�IBv"O�##"��F�XȲ�L��

��y�F���a�.)c�BQ� ��ybj�0�����d).߄aW/��y���)���Eb�:�Hu+&���y��~���w݃b)ƴrE�� �y2Iڰci��FK 
@����NV��yB��[�2A'��p�x��5�H��yBņ:[�6�3�ª[�28)��y�NrHvq�Ec��K��d87�yB�M+Z���Y���CBB��Ђ�y2fҵ~�� #փ
:����E�Z��y�r)��ɱ+����i��>�yb�� -����$��s@�B��yR�۹ �\��"GѸg��ͲS���yr��L�~�;��
c���w���y�1ezB�+@� �&��y����>CvhR�j�)���vk��y��T�a��d��cΆX5F<� ,ż�yB�1z�b}�G��Mc>�k�m��y�O\O�j9�LL�=+��
����yr�ΰ7ia3p%�MD�$�y�H �N��@�"�U@����T&�y"�;;�8y��N�$HĎ�À���y���I�FP)���9w�\� `I8�y�G�R�Ʃ#⣇5Z�ʴ���S*�yN��X��� �Q�~��]rrG���y��O�K{� ��|e�!8c���y�/?<$��痩o��P�IW��y��Q}�Mx"H$iU�B��3�yҧ?,%*,U�d��KB��y�O�>Sa�E:�Gg��ASkҋ�y�+۱J��%R�ː�#~Ip�A��yR��-�!��C�<}Fm�! ³�y�i�1oV%Ô�ϢK�;&���y�j�<Wt� 0�ޫ�����;�y�ɁB�(�G��
X*���C,M1�y¯̤X�p����L%V���/��y2����س��,O{���IZ��y¨�Q\(p{���CE���1�yBfݷ4��tJ$�C	"��q�X��y��^=��aÜ�:�EZQ&A8�yb�V�N��؂Bl&/�y+��	�ybc�}�ajr#5@����X�y�F�h�L�p��Z4K�Z��Pyb�ٗF�� p�� ��(9`E[�<Q��Ȑ�ţ�f�m�����G�W�<��j�E��)m o�8������yª�%�n�2�o�w��T�6픵�y2 �[�8����ے�\�"�y���<��aaF\�P��5����y" �M���`T��k�,�y�A��7Â �@��8Z&�$*"�ń�y���wl��S�S��qA@�y��,����F����RQ�ɩ�y�lJ�qp@A��9��5�y��¢I��ȄY�Hܾ�I����y�E���qqv$�i�2ݙ�����y
� �\�CDӉPP:M@�L�>.p��"Or�A� Y���ɁJ�1i�H��"O��	���8�z}�1�I*��`"O�$�D
��P#�a��j�#x��{p"O��,'t����V��+]RA��'��D9��Q4��-I�$��l�Ic�O���d��wȞ��Z*����Ag<g8����<a�}�e���I5�@b��.^J�H�ȓ��*��̀N�j�f�2���ȓ,�N�;$�
V����A���tbz���Y�`]SA���m
�.^�F����ȓ|C�ȸ�Ŝ]Fz��Ӓ}�R�ȓ�tM�"^2i�rz�e��p�t��|o��c��-)�|@֧��"��$���	�y��`� �(S��Ұ���1�jC�.Ն�9G�\�-��lҡZ�~B�	87Ѯ��QR,h�����?�TB�I(F�$���c�4��4��?T<B䉴)L�t��-K�kwDT�7ˁ�t�B�	��]���!_�jCFb��C��-2Z�P���6V[V,�6Qِ�t��	;dwM���(:&H����{��C�&Il>�	���Hi0YؔLV��:C�B���cCB���O C䉶>��:��F���5���� 8��B��q���2+�4�`=�������B䉛�x���MШc�$�Xe�1�B�	0�tiQ�mЛ2S����M�1Ң�=	�<|y�,�!>����n�%< z��ȓj��(�̪C%�xJW�6�~4F{��'����NQ/ ����(X'I/H �	�'��!�cTq��b��I;ڱ��'"���n�/N�N�!C֫E$���'Q��:��m�����㙑@�h�a�'��К�JH5��B2E�;��5(+O&���S�L�$����%p;�1�F��h=��Q7o,D��R�c�i�	�Q�������,D���G�/TS���G���@	���$D��{ԈD�ER�ݹ�/87�\�!�!D�D��f��/
����� b4�!��>D�l� #,��H:��=m�>�R��=D��!�Ȇ�~��!(㮔�/���p�!�O����OP���<�O�1O~mS�ˉ�gU�@:7L�U�Akb"Oda�΅4d-��������n���"O�6�ݮ4m`5ʴ�19|�f"O��`G�ݷ��=���v�S�"O\({�)@¾l���ɫ2�\1I�"Op�Q��vP|�b�@�$��(���'��Y,[I��)��Q�� ��+��Iy��(��i��*G��)��+� (��t�f�|��'s�� �ռU(�n�KU씐�'�B�V�[�`��E���-�4Q0�'�Y�D�٫*Z����"�l�K�'��� e��
e�MZ�DȖ#(T`��O�e����w�,�0��	D�S��'U�����cִ�X�j�`���Ȧ%1�D!�SܧL��ҕ���>;R� D��4W�Z`��pr��/\U9J岧�ވ?����w�Z��MK�8"0Zw��7�����r*�Yj��v_��a�dΜU�TQ�ȓj�T�Ҳ��?%θ�Y'"P  i���m�'�&a`�� �
v��
3D��pY!���)�D&-)��m��A�ӽ �����A�'�d�� 8�՛��m����
��� $Ļ�F�9@��s�/�9z�b���"O�r�B-�ⵒ#h\6]�>�H�"O�x��r�~xqQ��!w��k�"O�q���c�h=ʷ��������'�1OV�+^�G7ĝ˷��9��aۗ"O��T��1i0���ҥy�:��7"O�$+'�̪�.���䇣T8�t��"O>���ΨK瘥z$���I(2��E"O�h�C�r+�up	�� 5�m"O�Y�Vnݬ?}�!*r9��<JB"OV�iQJ�<Z@dH�H�&R�s��'���BC����Q���Bg��Ya� !D�������QT��J��DḰ�7L)D��i ��bj�<3!ݤ[�i� �%D�Z�Iܪ���i�,�'~>�c�"D�,�2��"q��I� U7:x.�1��&D�HE��:>G����g�]o�h�#%D��Ub܉|��s�-Y� �(� �'|O
c�x����\�R�cʼ,a����d&D��`�85�쁱���X$`��&D�ȫ&OL�Y-�������`Px�4B%D�H���/=�)��L�$?�T�TM5D���g�
���FI:(>��9C4D���g��GɒhIEoG^�(�3D�lJ
V�OZ �Y'�y�S�)=D�BWo�!N.�pV�, X5I$�:D���SC��C$â
 �A��Oh�D��I�W��Up�a��$@`�1Jj!�䄆a<�8�Q�.�l@�[(8F!�d�!Z֐L��h�Wl�1�Q.!�d},���*�Gh�Ҁ���{!�Z�&y5[�`�� *(x���.�!�d�(�r��d@�+��cÚ�}�!��%�L�c`K3F-ے�- �r�|rQ�"~2�'p���F�2��ݴ�y����.q�2�xt&�5Lc��7��%���E�w��sJF0���ȓ	�@y��))Z�vXd���4�]��HZ�Sa�68�����ߧUJ��?a����'���!�	Rc�+V����E'��0C�I1�����,�H����"b����F{J?]S�ʺ\D��3ǁ
 ���+�2��U���SbR�jB�]a6�Pqo�+>�B�:�2P��&�я,F�B�	#lfF��qm�r�Iq�U�C�ɨ5�L����E.a�U�s�ԱK�J�=���?���Dִ�T=���V�lwF-@�c&��?9����O�@�Ku�L�<b��*@ĜK�5
�'ۮH����4� ����=cJxJ���hO?ٹU�H
n�DY�Gy��\a�lPT�<�TfO����駬� �܌�gDVI�<1��E�)Z�	�����XZ�<!s	�]_0�i���� 8R�(U#[Sx���'��	�g�/`@h�b��-U�0����hO����)�Ʃ�6,֐H�z�Ӱτ�2�P�'9���!��~6`K�̴2|�}*��$>�4��⬊ �*�C#ʄ�!Wb�P�"O�u�#�'���:�@l�<��"O��AAHF�Y��� �� ,�0"O�h����t��Ѧ͆!g~���'������cHP�ĵ���ѺU��yr��?�֜I�.(s��@+��W$�$˓�0?�� �&y>�i8�聙�dԚ"hGj�<�.[S��1L��L�q*�t�'�ax
� ����+D��0�S��$u�Z�`"O���R�&��+P!�6�b "O��{U�X(56y�BKE�z�2="O��kP 
p~tzP
���hq��"O`<��M\�,��3k�1n yg"O2��C��+�5�e�Z�~r�y�"Oq�S�ٖ8,��P�F��cE���"O:���x�%cFۨj	@�"�"OAĥ��@���܍-M���P"OL�AƤ�+q\�*p���2<�-1""O\5�u����$*�¡��'8!�$
n��Ȁ�I5)5�|2�ǂ�.�!���E	p0��� G-\U��%�U��c��(��@�FΟ�q���1]]B�˃"O���`̑&ﬀ��`�&�4rQ"O`��1S���Cu�[=�01�"O�(@����� t)�8$����S"O@fc��A�޸���
+l��"O��j K�FK�%[��>�1E"O�ܣ��0h�
B��|�2��D2�S��:�<Y��5>�li�@��G!�C!~�~�pP�Ա����)�O!�Us�)Ӆ�Ip|t)ؖ*�<y!�d�4XkT�`Ū_�z̩��.^k!��G�D����F^��=��fF�T!��t����&ȝ�'l�����p	!�+$$8XPD�_�θ��k�>�!��N�oΘ���ិc|V�A@��[�	\��t���I�h%�q���A�F��[B!�D�" +�m��bA�!t��
�Xq,!�$Z<�J�P`,+'n 8��ϐPD!���h�@��i�������(!��@,q1D��bm@R�HZ�&�G!�Ļ'�r�iź3H��B��ޠD#!�$�>���u�N�E`�a��] # !�+݀����V)D3�@s��{r!�ē�n)|eh�?M�����\=W�!�$̯61�t,�&o*�l{6 B�g�!򤙰?�t-*�#ٽ)�쥁�N�9~!�$GRB��(Eʂ�Y�@�ҢM�3h!�Ĉ�q�LY�R^Po�U6f�-.I!��ءT�"a���(CU����Ő{*!��>u�xR�!F5Zya���w!�����H��6�PUQ"��	�!��5*E��v�l��-h�!��غN�l9
�e�#��	��X+d��)�'|���C�c��b�VTA����3��Iy�'"h��Ȕ�P�l�B�0)j?9�Ȕ��*Z� p�A��~�Pϓ�O.���G)7.jpsF�ӱ�t�B"O~���hؚNW,��VET4~J<�"O6A�@蜈(Դ�S��Q�In\i1"OL��r�AO�D��R��
�4yҴ"Oظ��N��X��]2Dȇ=&����D"O��
���������"g�Q�r�'�b�|��T8�vY���>T"��7lӋ ��{��	(7�h\�Ce�
\9��Ԓ)�!�ˀA���#��F�z��%7h!���FL�!R��l@@C�bɣ)g!�V�%�ޥ�F�@u9��k"o!򄑷	�)!p��+�.��B-�gY!�d@0%�6M"��48+)�r뙊WF�y��	�!m������4yvA0&N�R@���d$?a`�a�b�YrGP+��$�NQS�<�  �
�)V�%����uj�ڒ ��"O´PR��$:�	���>ƴ8S%"O����Z�)R�͙�r�~="Ot��2A�<k���	����"O���Ӗ�0��CȣS�vZ�'��d��A�j�3�ύ0��}BfɌ��!򄂻\�YA���"U��\7!򄚡,\*���K�`b��Ę;�!򤑷�셉兏�/`t�Jv�ӚV�!�Y�k�J���[	���qu��2O��)�'V��Dc`�A�1����&*�/xj�5��'�m:#m�1�9;V��)v�np��'[���5�ٱ'Nx��&X�vּiXL>YI>9��	I+x��c���	D͋<L!�d�U�� �&���*���t
V�>!��B�)���A��ԫ �
�����y!�$�'%�p�eZ��؀a��s�!����,���Y�EB�8��ף0�!��-Dd袣�M�v�Q���9�!���is�XgI #&����c�mi!�$�>gPNp�iɣX�H���b���!�V.J*q�G�)5�TE9��S0#�!�D�`���Bt	�(X�����ХP�!��N�`8ੈ�C]�:��� ts���'��'z�)�3}R�:-E�-{���P4���fN�y�� �>P(�ͼN���6�L��yB�F�'����W�C�0Z��I5�yR�Ճ;\�����R�]��璟�y�Y cY"`IHZF`��3�"�=�yr��	��	d��7`�5�t�Ȗ�?��4�X#<��=MT��	�O,)�TiiDOe�<��$Y0ѹ��?~1�Pi��|�<AǍ�&�j��VL�lˊ9�4Yx�<1�G�N�xB�G<�rH2�v�<1Īϻm�6U���;�&���ȗs�<9�h�{wXUh�ņ�j@����p�<��.سi��#L�(��`"N�C�<�e�Yu��	"1
0i`����<��J*d�sE78���+�Et�<2�A�w��0A4)�2)�Z�͒q�<Y!�KƊ$�g�D�n*����Pt�<1��d��u�1c�/qR !���FW�<�p����j�%���9;�J�S�<�FEH8>�Tz��q%F`S�%QL�<�gz��kT�^s��`��Jx��Dx2��z�Ip` Ֆ[� �*adߒ�y ؄=�̝��I��g�d ����4�yB�=7�=z�LO�[wz�Y`�;�y��C'�Re�0��:J��L9WG�!�y҇��L {�E�mL��$�y�V6fr���N�f
(Y�!�+�y���?���"� ��^Ī�Q��ٿ�yb�_/�̬cE��6Vm�L�쒚�y�W�$=|� ���4f���@C�,�y"��ub��+���`|�Љ�T�yҧ)�,b�"�V��]���P>�y�솫PA�4�vS>���q��"�y��<^|j�@Qk� ,L�� P�y��\>�9 foX���(C�lJ��y�ӴM��i#E��8G<�Ӓ�ݣ�y�OL�Z���j���=c(��_��hO���N� ��)q��?v&E9b�!�TB��1w�܋$�\��abJ�w�!�Dʍ+�z��79���k1�Ӊ�!�� ���#�W�N#�����Zo�9B�|��)�ӌzV���FI��Ȭ���13,B�	�^���ū�� �+���*��C�I�n���eۗmnr��F)�D�lB�I������k�14�Zaƕ�R@B�Io����+	@�A��g�6�C�B��YHc'S=*T�%B���C䉶\��Uj�C�c�����Ϙ�c5���?y���IҎ-��rUDڔL(�䤉1O�!��D�EW 00�*�{~�@"�6"y!�@�a�V�PS���l!c��ԏ!!�[j��B��:A�D �c
y�!�����*�!D ��t��#��!�$̂T�T���I����6oX!�ԥSs�ԃ����	0�'A�$�!��@Y��1�S'��rc��3���'�!�d�P�h�P�/z^��h5L /�!��	�wX"���L	�Q��YY�*M
!�!���#���TLLO딬�1CS�
$!��ʅ�T�c�b�]C��``�4{!�d�	>��4)]ju�p�;y!�$x2�ma�$������kڂr!�䊈�nI�L����*9��'���'��4u��.cZ�3%3Lو�
�'���C�ůPb&�J&ER��I�'�P��D�Q?"�V0pA�5��XJ�'�J�����t̡���&v��0�' l�Pa�о�Ƞ��&ę6v��'{\��H�&?`X��֍B˾�L>a����� .����ˌ9n�-2A�N�>��O���N�7� ��'EW�B��kSR�!��!)�<��O�~H`c���+�!�D�D��}j��ė}/j 8�
��	U�����D7���i�Ƅ�%�&�1 ?D���֊�B�B��؉R���9�=D�0S4��^(���SȔ�%n=��5D����@C�,,AR�A�A�z���-2�� �O����<p8ZfeD:*8dje"O��PC��T{B�䎉�;'H�@"O�h`��oϦ�B���f*�rV"O�:BOC>�&��uoކ��D��"O�H`�
D
�����s5f��"O��a��C�}���4]>r(�d"O<�+���!gFbG�hz� �Z���'R�'E�� c{�$}��� p���'R��T,V"�����@�&��Y �'g�郀h[0_�,z'*K��>��'<�k��%
�ҡ�uNY����'�X���t�#��ݦz����'�l�"Oȓ��P�'���'Zt���J��N�Ќ���O/���N>����0=�b ,ص���/: \����V�<a���SPD�	�Ι�����Q�In�Dz K	~nd��oS�zy ��C;D�,��ǍC�~��$UR��c� 5D���.ck��TG͢8�p�
�B4D��d����0����w[�tk�6D�,�Ԯ]4K�<m�E�����{��4�O ��)2�kĵ	����ǉv�T�ȓX8�Q��_�����D�L|:���eѼZ$�P>\�8��"݃f��@��(�6��6h#.]�(ֿk����� �0M"�H�vD2��-ΐj4��0.����^8ef� )����l���S�? ����ɷV|�����ȍO�$D��"O.��J
;F:�`ß�M��B�"O�e1�
�Ƙq�F����{�]�H����*:��3�ڀ#ʹ|�fj��\�C�ɠ6h^��G�����T+q��,fxC�+;�`e:�Ɩ�@�2V-aZC�əixEKW��TވD���0�4C�I�5�,c7N�T�(eRդ��$�0C䉦��D�dZ�&����O�v��C�I*x����A$OA؜˶
��(���O�����Y1.CIC�<�,���L�J�!��Õ-��M��.�R�d<�:��'���ʷ�&���˘
:�h�
�'0D�ԡM�7�p��E#7H Q�
�'����G!D���!MZ4t�	Y	�'pZ�
��Pu;��0��(b�=��'��41fIەR?��H��]Lk�����'X�ݣtMC'{�h��f�4K�z���'=F�hu�Y�Z�&���MR�ҡ0�'�`l�qI�m2�N��H���r�'ꠣ�g�Re�1��T[�%Ӑ�y2�R�N�VI��^��n��e�Pyb �v��B�.��s���Ȑ��V�<�1@��D��9'%� K����P*�Q�IΟ8��I�K��er!�X�C2|�r*͐zڌB䉰
J½���6n�f<I���?r��C�I�&�����LHF��*��E�}�PB�ɖ)�$�k�8���	F��B�	%?�9�픙d:�9R�,H�'k�B�I$>\�%1�� g}�Q�@?f�^B�I�06^�AN[3(��qS�Q
z]LB䉌Wr�)��*Z;�ĭpt���s��C�e����K�<���3�N�F�C��ج�� �]�:�(��Č�WHRB�I$;L�D�BH�m� �Qd���C�I1GM�9rp�W�#Ti���{/�C�I14!�Eu��%Q@h�)PE�C��8;�P�Æʝ?��eT��GkxB�ɷ)���lB4?~���i��4�C䉷/� �%��\��M26�� �C�	:��*0�(;�;e�)�C�I%4Q� ۃٕx�T����yTtC��:H� ��FG�I�1��&]�LC�7̂t�!eC8R>8L�vݸC�C�	�iyh��'�@�&
�����2@Q�C��(->��[@K]�JS���6&�./?�C�&�%(`�B�`��.2E�C�>Z�ܥ��ā?�j%C��Y�X�C�$��A�t��~\{w��A��B�	��d�8��?R`�ī�v�O~�d1��O���8?!ĮZ�[H�Mu�_VU!�X�<��e�H��ˤ���#
M9�Z�<�  	IbA���(�����W�<!�@ړ��x��K;�rݚ�ƞQ�<A��mD$s�푼eB>$Ð�e�<��ˎ�zٶXz�E�,U�̈�!^�<w�X�1<td��Úh RU��Dqyb�'7��'ѐ!Z�ۘF�*|{AY$8J���')b)Ae��Hb(9��C��4y��'+Ľ����<A����W��m	�'�lxXA(��ex�E �����'=4	�̃3��
���sD�	�'oj��k�#S�i+Z8� ��l�a�2�ΣLEjhx� Z����S�? �As0�V�/�5)� I;���"O��Ӣ�\����2	� ��Qa"O��!�P*�Sb-R�D�TE��"O>M�ԦC�AԶ�jPl�<-��B�"O�����_+*��!�4��6M���Q"O��q�߲j���K��k�j���"O�� ��J� |�Ae�4>��t��"O6�
�聖'orPI�4���k�"O�x(���8#����F�k9
p[#"O��ÆCU)&��-����&
)H�P"O�}�7A��n�\��q�U	"����#"O�=A1HJ�GX���GX<^B@���"OZ��e�Q�V1�qFbܜ��"O�E�EY�0�Ȅ��ɕ���(�"O.���h�l��au�Sp��@�"Oni�VJ�'�r��TJ^��"�"O��T✘,�<QE��V��"O6��u�!��Iks�I"q`���"O�	��"F�t��RG)�-U��T�A"OZ�"B��5v���@��N�d"O��+]��=+��4t���2OP=#��D�;��G�S9��p�� D�x����xz�����^�K�$D�ș�� -L��Cg�+{F*��%�#D�t�"rDx����%`��0s!D�< b�h���	�IW�k����� D��`��B-3��,�FŁ�'�`r��2�O�}��5�1eޢO��(x��˔P�
���ID̓R���ECPa�4��0���J��Յȓ6?��h�͖.���C�Q���P�ȓ-�Na��L�7Vbrœ"�B�^ ��.�\�U�8f� ���e�<��ҋl.,�A쐴P��qe�6d���n��d�0��)�*2����"OV�Z���?P0l�u\�����d�O���O�K�G�9)�C"ĥ�U6�yhؗ�*ق�!�K��D��ʒ'�y�m�5^)ʓ �7NFp�'oV��yrN
�8��	�Ӥ�|��2͍<�y2�/@���b�䌁v�u���y�h	�\�ΰ�g.�q*���T�\���>����y�gM�(숛�E�/o���B�����?���D@^X˪��w�N���Y�	�y�@
6	�X�{|����\�y���^<*�:�-�
�f� ��y��L*�r�C�, �9��B<�yB�6?�"�˳�ef)�&��yl2`~̓�n�9�z��� Ɖ��>���y�C�Ib�ĉ�'k��R��,�yڤ6]���QM zp����W$
z!�D (�L�PW��,`�I6
XY�!���S�xf��&5X���0��S�!�$�p�����M8�}Q�*��@�!�d)Rj������L�C�A��!�
!{ �Q�ǻ>x^E�&
�"��I埴�	l�)ʧ>�41� ��gEI�4E�(y����lc�!hBL�g�N�)ՉQ�t��U�ȓA"��XRB/G����Յ`ꩆ�z����Ƕ9Üm*$c�9/��(��x4V(q�˓.J-��*t��/P�8��z\=	�H�GZ:��º��y�ȓ:X`�XU�O6R�d�zP��/؄�	ɟX��� ����dd,��c����0��;.Ÿ�OL��ƮR��l��L�5f�U���r�!�� f���T��ocS<$��e!�"O�� A�b|d�KPb#��� "O�HS���Nz|��!-H`�Kr"O�m�7�$N׀��B��S��ٺ"OXL�U�[*j���hK�r��Q���';�'��)��t�!���_�]�4Bș{�*t�
�'�t@`�cF�`��,	#*vb��
�'3PI�E�.}� ���p��ma�'Ԣ=���1<V�%��G�h=��)
�'u�b4#TFU
�K��q:��Y�'LV�:�I��A�6�h�Z���
�'�8�X�G�1;`V�["��F�  ��]bp�@�_l��OP�_jJ�ȓ,X�!Κ�Mf���V��2��L�ȓ@r�	�S.ء��U6K3XB,��RȲLp�I-�l=�S��vy���I)>�F�.Q��A`	]|�9�ȓ5BT�k�Fl$��B���+|��'���Y ��?�̬�4H�F�"�'�B�o:Tl�S�O��"����?��_2B=�P�J�0V���-]���ȓ`JtL��K�6y��O*���ȓ7Hr�y�gG�3b����B"fh&����<��Ia-b��k\4𞥆ȓ3�_+-�&��D��,�i��	�02��܏-B� w�x�ƅ�ȓS  �bR=t���s-�^��Q�����Im��#�	(�e��$I>�0�I&D���A�'�*�Ei��c4ցxQ!#D�$��mP���ds�/>7�����"D���Ig��C
ָ3������"D�,0���	C<�2J��HE� D� "#���.�^q#t�ͥ�BPI�� D�d[�%���` ����(��4��
>D���AfŔ%������v��x��l:D���d�'l`A*���"��(�"�8D��ԍV�
� ��A�K��BT��5D����d��ؘ��%�tD�0'B3D�@EK�P@�|�db�.4f,���2D����̠E"��{F�x�l/D�T1W�\�0�� q�˿X�!��;D���UځX���X$��-6|밪<D���5��Z�AZ,\�}�����;D�hag
W�u��	!�1��$�h8D��R�LM�sҰ+�@�xǾ�s /7D�x	��	�X�hDS$G�%%B���)2D��Ӡ��w;L��`I����Ջ.D����\# ��8��:!`V�*D��c� ��MD������{�ȩRA�(D��	�n�o?Vm�A� �R��� �&D��#%1u����#	�:?�IQ�N D�l�6��$� m�ԢǮU�Lqb3a<D�
��>dp%���E�bY��x5-9D�@BFI�%� 1� ��%Vi�V�<D����폚>r|�W�\DL��r6)>D��#��Hkx�H��<{<Xa�v�<�#��w��"�T;z2�m�wC�X�<��oĿ��𡒄P j㌵çhBX�<q ��D0FA��Ίp6�J�o�<�ff�) ���Zt.[�Mv���o�<�兞p�`Y�S�Ƒ�����N�C�<�I]3&�\�#�I��0(���x�<yv
,Y��qР^4~xr���IO�<��c�	\�9�oL+?Bn�˦��K�<� ��k��̊A@*}��i1ɮ(�2"Ox0���Q��9�g�§1UJX�C"O:���#U:P� � FT^@9"O0�����.������EO���W"O�qۇ�+6����	bj���"OP !��E�5�pdJ_�Hh� �'E�y"�d�9�8��Ai�^]Ys�9h�!�$ºd��%pE�Ȥu��d��gU�=�!�D�-#0Tx�gB5td\�g�L�!��;���f�+{V��bi͉m!�D�-_�ABu@�F��iݚ.�!�ԉ1
)��
+AlL�g��"�!�����8&�8<�IC23�.0���?����O@�h��������I���*P#ZP�ȓIm2`AqB�9��m���Ϧ'R|Ԇȓb	$X
à�oo����V�d4\A��l0�����I55i�ȇ�¸}�<�ȓ<*@a��Yx&(Pf�-a�H����q��c��{���uK�*Z��ȓ�<H�!�w�A� ���%�}�'a~b�Ô2�"՚ %,��iB��y��Q5C�&pc�F�>���kޙ�y�埒4��4Ka�_;�4a�@���yҍ�0fft��(K"6�F�2����y�\�i�����%+\L���W/�yb�VF�`��W�����"a+�y��2�\Aj#n�"�V�� ���yRH��!Pn��oE�.�c��y���,}���F])C������y"���#ɖ�𣖖i[~�B�yb`D*&'��ƃL���bJh	��E9�	�秏?@I�iO�ve���ȓRK^�q@(��|�l�֏�#�<�ȓ��T��GJ#A� Д@�I���ȓG�1c+@3zr�D��#��`�r݇ȓ�R��Q��$�N�" ���\���9���؅"1T�������	`�D|�ȓX��Aaaξ0�d�z�*	��U�����c3.�|x�
���.�<T��S�u�/�����[���+:Kb$�ȓ/;�T�WO�T|X���+~�D��Ox��htIҘq�R8��l�\M���w�,�	2��F%н:W�U_І��l%��ۉ,p�ĩW�^�=p��ȓu�$Y7��p�B<)gm
�0�ȓ#f0 �-��}| ����ǂ;�v��ȓ&A(����ɖ�@akb,ĉ'i�|��J��Ƥ]8p���r%]	M�"	�ȓ�~�Bċ=4�X��Ɔv b��ȓ`�9`�L\�Zc�䳧JΝ4J"ԇ�
� ��A˲G.�3P+�����ȓB3*��&��?,4H�7E ��tE��*)c��B�L����s��e�m��L���b獼Yf,���`ÕvN��ȓR*��dK&-������5<X �ȓ�q@fS G�ᒥK�O��ć�y.,7��BA�x*���4%�,��"���E��% ���"�_C)�Մ����d$T� �n0���Ih��ȓ����Ơ�OD��uJ��1�6̅ȓ�lЈwI���D$��L�L�������'� ;w��Y� īQ��t��'�z����V�� X����)����ȓr���B���q�(�CD&+2���S�? V�9g�[�\����͛&����!"O��{�g�$5�(�K��0Q�B��s"O:=p�h�0/�Tx&��a��@�"O�ib�$� 6�$��a��ẹ��"OR�P�hܥ}�Vm�
{����r"O�1�b��[��K\�dY"�r"O|��\t��ٺ��@8TO�{"O��B�
 fj.��GɌ�@p8�!"O�\2���x���>���"OR��G��*%j��A���4f=�%Ӷ"OL�����@�$�uې;�"O~�@qI;R��H��/�'��|��"O�)CC�*t��	$�K-R	�%"�"O����!Y��e��Ό2iL1��"O�� a�˂Z�(h�$EA�~l{�"O��[�#�`���Aݖ�tIc "O��:�	ֿT�V�3��?Dt�x�"O����,Yh*��A��63��!&"O�!��*Y'ʀ(��N$&+�i�"O��0�bɄFW@d*a�])d�`:`"O��(Q��J;`�)Wٌx|�(H"O��xt ;B$���)�v���"O�\`n��\,.-��u�Hx�"O^1XQ��={�ЁU��w�ȅ�#"O�H��ڍ'z��vL�)(��!K"OP�ZGk�n!��[嚩i�t,p$"O��׋]��}��d��c�*�B"O8�:_(�a	��/���h���!�*ELT��d��]?�&1D�!�< P��� ���:2�4(!��$\Q��(��ޙ��y��=0!��b��%���ˬJ��WBſLk!�Z
"ұ�a�Q�;�`�
�A�51G!�ڋP\	�w�[K�<��$��$BN!�dțez�tQ�%Ҕ�<���H�#�!�J.VS@!@�X4.tk��ED�!�D��iN}qA%�<"�I�F�Q�ky!�dS�i�)���CX���R�!�JZZ��3� T�~�L�iW��!�D�I�VlȢn�#��0+�Bҿ{	!�
��p��T�2`�$�S�v�!򤝞#�V�K�N�t�R�B#;�!�#1j>mS�.\�*�nЛ'.!N�!���@QI�!�%/�~�فl��!�*���B!o��<�4i��V4J�!�d�  Z�T�]�V"�T��"ڗ5!�D��(f<cE˘��Dc�J�JN!��<-f��ӥZ4x���d�A�0;!�D��fUʦ���H���^D/!�$�1d]>UD�~K���t�£f%!�W��9���G! 61g��9�!�$�#�Fd���ȗĢl�e�GB!���2�d���Q�|����)�Z��'��M��"%ua�	d�""��	�'K��JÌ�ahp��K�!4j�'\\a'���B���B��>L:�',8�$�P� 
��s�ET.	�-H�'�Ҭ�3�F;B#�4	�͋}46,`�'����JD2=N�ـ��?u!~9�
�'
^�ccIuj̍��>n2�	R
�'^�T�2�СfC\�ㆊ�q(��:
�'G�A٥�Z�'�@�� �7R]�	�'�ѳ�l�;ߺP�ŧ_���٨	�'[M:�ʁx���: ^��.Ȁ��� T���b��:�]6���q�L��"O����|9eڳ���U��	�p"OH`��$���U��D�"ٞ�!�"O�%k�o	f��hC=_���9�"O�iB&/��V� ���F3=���x�"O��Q�O�I-VA�`����0U"O��P���7O֞n��B�"O`Eҳ�\E��l�q ]�P	ѷ"O��@�D�%���u�ӡ��%V"O������H}b$�!�\.4��QZ0"O�ASσ9_X$�U�]�s�bL��"O��XC�D��`끱����"O~���M�PcV��u���+�"OX0�0V�)H�E���7ԍӣ"O$���v!���1���Q̴g"O.��Z�6I��`�G�CFte��"O�P�w�x)t*]r*R��"O�x9�"ǱO�UH1��	����"O0ɋ�׽k :����!
ڀ\��"O�Lj�J�mq�e�U�D"ZŨ��1"O"�`���xb� "��d�V"O�Xp4F���}����V�~Kf"O6��3Kٮ*+p i7��p��ı"OrX�5��d� ,�U������6"O��h�L +�n�JiܚT�A��"O��f!L2Y I����<W�� � "O��A�O$O�%��><\��"O�<C��%zp�e�`��=>.<Q�"O�XR �82�|�IW���Re"O^ ��%�']?4-:�g�=8�� "O���H7\�����3�T�kU"O�V#S<i���q
W����"OT�pRO�#l��G9N���+5"OdW��3lK��Y��N%b���K�"O�0���I/��9���u�4�D"O���qY�1$Ȅ�E��3�Fh��"O��Wd�7\|N�	t� �13"O8� +
������%k����B"O�x�V� 2f�F��V�µ#v��E"OX���R�((l��K�Q��!�"O��駉ѐ���K�%�:oU|,+C"O(,� Ďu��H��(Tx��"O�-⋁�.y聛�@�V9R�"O��c�E�*��	J�,s�j�"Oj8Q�F�hit�F�B����V"O�`�e�?U$ȡYl5�"O�t����RLZ)b0��"��(�"O�ɻe!?!�L0�
�0d~$u"O�p��B@�m.��rGCG4O^��"O�B��?`K��d ��3-䑩b"O:0a�j�13肴�M��S%ڵ�"O`x�D��:v���%ؑjz�"Oj�B��K 
�Z̋4�G�XX�"O� ��A�p��!a��8 ���`"O@@R�@��1ɬ��dſ]��"OjRLG�v��A*d/?U��p"O�Hp�!�!-̥����&8���b"OF�ɶ�@�炌����X*N!��"Ob}��ˉ�:n�-�Cۗ��q$"O!�鎀H��P�M��
�!"O13�c8�D�21�@�rq,��4�'B�'������ƞ.b�y"��%��I�	�'DpLH�C���!E�F�TX�'3Ψ��!��aʨ�P"*8E�҄��2�)�� �$�D�*?��pHE	t��2�"O\�S!��8�ع��bM�%d̽۴�	S}���++y�4y�M��W�P��冔�zQ�B�I8\*.�j���_���c*E=-�O�=�~�dD(2��AC��L<G�5 ��G�<��I*)��h��:+!j�C���M̓}��X%����$f�@q@�WgEv��$��7O\�3W�F*�,J$���"�"�OΣ=E����.(�(q�mK,��XJ�K����'��Ix��u� Z&���k6OO��ଳ����x�ED�j 6�`�Aݻv\�&��,[���E�d�ą���`KX��`�ꔴ�y�'m7��b�C�=u��W�W�y2�+I,�d��l� ���Aș��y�b�K�^u+C��Sl	��/U�yb�� <�e�#�Y�8�|1��d��y2	�9Vu�\�1 Ϟ2��PP�"���y2�޵zE0M�u��\*�1�Β��hO���z�'��|k�$U,3����.��ybC�>�,��!7�Y�`�*6�C�	2Y�6��
9�PY�,#�j��D5?A��S���Mԧբ�۠�Q}R�'P��� H�]yRxҔ�kڕ��{��)�	5$�.�L���!��lѯ`z!�DJ=�"�x�O�+rזa����0Mk� F:O��=�Gb��Ua�`4�\�S����xb5O�-���F"6-�0 Ϯ]���w.���E{��I7V�����z"���yB��P�"m�g_�0��)�)���0>ّm��qB�0��F�:n�P1��@w�<1�@�4+U�@�e/4@	FY0�v�<���ҕG�����Co"��+��u���?a�L)I��x�6년G�
�es8��&�+!�Γ&�؉�f��Yz���s/7D��F�h��P�(\n#��9c�3D�Ȱ�L�;`e�?w���Q�,D�l��O�?\� I�v�[�i�lຕ��&�hO?��o���'�k�[�̞���#�}2�Fox��a�ڷO��*�L$x��~��'&��Xf��2%���U�-U_�x�'�*��C����
՛nL�Sҁ��'�,�`�Ń�O�b�6a��R�#��d4�^�v ��p� /i;ԙ����<�O>!)O?e�gc_� b1��%U	{O�(�C麟�E{�/�m�z��aͬ9��㥌 ����<��?s�|�#-w8 ��C�E����O`6�!�S�'9��l2���
h(�����68A���IGy�DY�a�	��㊌B>��iF&֏�yBɘ*58r��A�@q��h��xbLM"I׆���(����glH�V4ZB�I�g�$	#� 
(����/H�B����mQҧ[?(�p�Ѳ$k����'�l<+�es�޼BҬH)h�.ur���"�	�cu� B���gՈp��B"A�B�	
�t4[�*��~�xep���=�*��
�'�`���ǈ����a���*&@xT1��$��$�'��	�`���.U�(�CI��Y\C�ɽ���p�J
�z8U��IYY�\O�ʓ��S�r;�d)g/bԬ�	�V�q��)hH�� &E%�$�H�<��ԒR	�P���O[���k��l�E��_���R���4&4����(|����%��0�8Y�"b]�:�mF{��O�䁣�?8,$�FLGX��yO>y�����,6s��3B�Z���̡�-׀'�2�)⧹� L(B'͖�#��쀷%ܦ:ø�*�E4�Sܧ����O��o�"����Rj;jͨ��T����	�G��9�$I�cUx�����'��	G����3���՘��F�Z����U�!D�dq0C�G&ȳ�i�"2��
��=D��*�eI�(|�)���.p�\���;D�� ��Q�!w��T`Ú}㬌���7D�����,-d�0��B�L�B���*D���u�C�@p*㦝��B�3�;D����!� $t���rC7cj�fg:?	�i��E���H�oP2�C� �g��P��W�4��S�E�ϒ�[�S=<r ��8�.�!��V�U�t8���P0�D}b�yP����X?�L�(�NR�B�	�tm�U�4��-l �Q����	�pB�>S����"� �ub�d�0T��B��@�@=�%C�a��@b�X	��B䉊#�L�!B��n�M��/T&3s�C�%+�: XE }��%3� U�m��C�(R�\�st�O�	�� �N��z��'F� r�/��Lcح�-ǟ.*���'њ���I�*t���d��	��p��'Ge��'X�|(d!"��ǧ���'���(a
�M�~m{#�[Մ����(�X])�"��P�2؁��x5�<�ȓ-.��;F�����<Fw�"�_�Oj��� Ig���yv�ڝB�:l��'9��Z�aA K���".�8���
�y��'�`Q��B1*�fT@���[\޴0�'�B�׮�0���1٪K������x�;'s�JB�РNs6�34V;�ē�O\���%=e �sG�3w�8=vG�Z����P��?	�j�([^^�2�$�#
N A��AB\�<Q���7T���	x��I�" b�<a���y� bv�\hX�Ñ[y�'����Ӎ�<m��b�7��(�*O
�=�O�	�=��G�I��a�QL�jrC�N�3�-��7���C�<RzO�����F�p�b�֍w�����
�1?��r9Or����O�=SD��LH��� �"O��@�̐�x,^��t��"e��Ij�OкU�blF=8�*��J�	�l�:	�'����G�<Hv1��$ƻ���@(O�=E�O�:���RLۈ)��!S��͓�y�(G*~�$q٦�$��JeG��y�j /h��P5`H3�Q�7Y��<����sJ������*��AEm�en!���_�� �	�|JK�"HH�'Vў��-}�"�y�@xH��{��}��΢�y��!i��@P&anr0K�yr#Y_��9�^�M�����	�y"��9�J�s�
0Mѵ�M�'&�Q�b�-��"����j!��'Aj��H�ETf� G` ��T1�'�j����f�j1"�әu<��'� ��W*�,(H�Ԡ��ۅu��e;�'!Byh�Dǔ~?�1��i�v�q�'?���f��m��Q� ��.[��	�'��У��?>x����$�,!@�����6��9���C;�d���MZ�/K�x:"O��4���N��Y5�w!4�*�"O��%G�4FF���>��G"O@��h�:h��Q�JM2�6�k5"O�a�3�-s;�L����(83e"O� � Tc� f���� �!|捐�"O� 3�Q1�e� ��S���"O)y�$ۋ����T�݄L$��D"ON�	����(|b8�'#+`�𑈆"O<0�d��|cd��%B!����P"O� p7����-�d�ن�2�"OtyRv���`�xq��P��Fl��"O�t�tHϊf,��Z�#��}�ε	�"O����E�&rY����O;�1�a"O�ݙf�B�{y�!ˤ�%*)^u3�"O���R�O��l
�*j�= "OQ'���b��ل"� )�%"O8Q�2�6�|l���2nl�U"OH��E"���^ !�)��/���!�"O*� �] bv��R�A <��Ig"O�9ktH^��4a�m�h^\�B�"OJ-u�],/}����ʊ�K�<��"O>P�D��j�5G[$�H�"O�����=g��m*��A�"O��Yp/ �`�h����/�D���"O�Qiw�!t�M�u.�x-���"Oh�G����qp.J-$�H"O(� �RK���
$g����h7"O�4KS	ˡ@HthY��$�tIQ"O���h�&WfЉ@�g�M�2�I�"Oƴ����%{��Ou�"�"O��[�A,Cd`�;4%��ck<%Y!"OJ��W��?(X�����R^"O�	���O$C@��2Q�B0S�T�{s"OB%�`��:5��,u~dSW"O�X�DlKr��h{���a���"O�LC@"ð&�R�����I��"O���	�>?Ph�7I�.us��=g�^���'<�8�BJ�>ZءB��F#��r	�'��MÀ,E�f�2�`u��A)���'�:t[ψ"��581�͊?x���'���H�E,��!��_'+�P`�
�'?�Dq��R�{Xн��!E�A@
�'�zف���3a�x�%���2	�'G��'g�R(�@�r��e��'˂񐁂�:U" �8b�	;ܚQ�
�'}V`�`�չ`�<|��L&?��<�	�'mt`��K^��pR���*c�4�'��$�@�P�J���S���v��l)�'[��z��l�Zd�b)�cC�c�'���Y� �y@�U��J�K���0�'����CH�!�t�7�)��(	�'?F�� ��$�Z=�
 xT��'���E����v�P6��'> ���원= �[f$�02�b�'���pF5E&,y�bޒ}k�}#�'�PI�#V�g���"b��f�D��'h`����S�A�JS�])�8��'��UQ��9%�"Ā��ʸD:�2�'��dk!�
C�P��\�zg�:�'8f�¤��y�����w��� �'��XJB`$���l�4y��@�'��[���"�0t)��#`Pi��''��`&��N*��u��c�yJ�'w��!"k���x%��
�X�#
�'��H+g+@�~R���4bF��d	�'����5��/o-�)C��N	�@}A	�'���Ճ�1f��
\k��x�	�'@sO_�G,v��qÉ*d�
T���� V�x�A��N�)µb�MĊ}��"O$�Ti�:TԽ�'���T�kr"Oh1Z�@�c����%_�E[�<At"O �C���-���@���`8��s�"O��9��M�[1iph�w�USU��j���C8���!�O�-�z%��&^i��Qm$�O|��7d��y��$@�A	��ĩ2��І���yr��P��HIG&��3&$��*O��(O�����Q�ш��<�F+Ћe�4�0��$��}�"O,��ኁ$"�x����E�5��h����dB���OH�Ӱn��4D�ԑ!�ǹ@_~9A4"Oܨcr�ҟq6���_L!l���O���!OT.�0>��HF�.�!��SN����B[8�0�w �	o��K�'=��7�51*Y)tO-�!�dͺm�ک3�Θ<"Dpu�� �-wz�����]v�O�҉��9O��Q����qW��	�'P蠨G�M�	�,���Ԩ`��}�
�'�X�E��=w��<ˁ�؋a҂e��{�,�i�#;��L� �B���-�#>���K��b�!�d^w�l����)h���W�	7V��P�H+7/ ���S��ě+h�kD�;!��:�%��V��:(��y��ݠu�Ѩe��!��p*�iZro�	�O~i�4d51�Р3$ >��'��n2?��,�W(L*v��Y@#�4Z�!�$3<쪐�0	�z!��g�+I��%� �%�6� K�#{�'K�y:��ih��{��@�I1��ȯ8��T��-���u�4Cz�'v H�1�^�k���G%(ƴ��O~�h�n֦M7&Q��`�
qhN� 7cQӏ��j-�'l� ��F� 1�ݦO��'1��:�̗���0ᡭ_T����P�L�s*}�$O,-�pK�M��0���L�ƝJ�'�3���3���[u*N�`p�3�I�Y��ݼ˲�ȁ3�,��1/��S�T���_<��	ȃyb&e��CP�o\l����J'�Eɇf\25�f%����I��p �nڸg:�㶣T$��2�K*�����7�$<	 ���
�$�j��L�+�F�
����M̲�a}y�U�+O�(�Ҍ��5T�f-f��� z�+�L��	��)}Bn���;�|�O��	Yi�4�!�.;d�\E�"g�0����K�B�dN�	eIgl$��O��)%B���AC���7g"��x *��3B< wE�+@������xP�JQ%h��&�Bg0A�"��$MK�k��m��d��ɈB��-�%�'��Pc��F�o��KE�
�ݴj���Ї���!P�	�\�&с�(��{��Q���-��s�Y�"���G�� ذ��(��4��e4ʓI\NM�r 8�H� 9X"���ћ O�QQ<aPc$�'G��9�	?�TYueS7D�'L��� �'K(���w�>D��5!�$Pˤ��R)��qѫ�=w�A#�Bu�ԟ�U��5�y��:@����8p�RVeX9M@z4��Wk���Q�fR����ŢAL�B�'8r#=�c�Z�a��	��W ���m��<	��Jer`1�������eph-�� �jږᐣo[g]���'��E����$Z#@�I%�nzd�q�I�'�1J�C1*��-�7b��ZV@�q�ꍍ(�ܴ�p,C��T|�y�a�#�R0q򋋪=N�������q̻M��q0���6W��}�@d�V12lDx򊆇�&���Eu���4�	�	���BA�� ���X�5��T� j]�B<0���I�Mq�	�
���>��$�i}�0Q�h��+�x\�X�<�΀��'��.��B,Ge��O'/q ���N�������3�n����;��Iե.7�0ï�X��k� �0K�@m���1���D�"�]U:��(@���Y)��	b�p��i�C�	 r��b�����U&/�a��ce�x	T�
 w��D��N�(�@�A�t�cO�9K�����(��X�cKA�X}6�aQ��`����"]sɒU"V&�7�I
vr�+�I�~lVȀ"�Fb���PWg��a���ٷ6�JU��Ɂ��Ds���Kt5�4�I�D����f�U=�O�2y�m$0l��4a�*a�NR�W�;t�J�C�IΠ�!�p�N�:|���	�O ];�K)VܠXѣ�a.2�(R5���Z��
���	��B�
4-�L��U\���ך^?���v��1E#�Tۣ��@dz���#\�n�|C$�O*2�ψO�I�eԜjB����ѝjC\�J��O�L��?��D�ȹf��9-tɁfd���d�=@��D��D�(qbZM�����a}�G!a)�)��#�H��O�}hHy�0A�	Whv�'�Ԅ���3���@��	��	�f!V�љOo��81�%�t��Q��S�Q���*ִ�!�c����Q�6(DI���,m���h&����'�L)�q�Y��'.E2o�6�� /��r۾�Ja�q���h��=��8˸��4�#�I
Zۺ�x�I�"W}| F`@�3s�plڗ�(y;$�N� ��{R�D���p�&�n��%a�~��Nh�<!Dz©�^hjy������ ц��h��vAH�Zp��'3.�2a�H�<Y -��6fː`�8N�@
C��p�2������6//ޢ}"�	�'Z7|����R���EF�'Z�MXU�f�O����!Z����K�n*;g�@�д�ś>&�>�W)J�(�n庲��T}H;%��|����"	�n�S��?��/�<�8"��K� ����[���w�Ah�a�1�'�LT�B��5�$)�D���!h����'W��W�Ie�'M"�(�-��d���		X���u]
� %Km����V*�&�I�G�.P�� �g6͸�^�Lb�Dy�G��ūP�!rj�H�gL�OX�`�L:1�@B�	%�*��e�/�p����,z�@�pR?:_4��J����Ouꕂ9+*i1�$E}�t�D�'|��u@$��Dm���x�A�ė^C~�ϓI�B����/�O�1��ý]�r�BĜ*=�!��"O�M�#�X	�&�P�'��c��d�4"O�]sdH
;��uCf��w� X�"O� x��A(a��50G8\����p"O���2Nڜ߬x�¨�����$�i\�M�� ,v���Ki� ���(Q�ن�>�̊��4x$@���>��P2��L�	sL)��I�2ЁA(#�PR�J�B,���$��A"��#�<�r�R^L�D�B/TZS�t�f�}�<��l�|$���l�
6W<A�n�`?�IN�e�T�����#w�h��)�+��qUJ�c>�]�ec�x@!���Fj�0��ꁎ:\�9��Y�K��+Ħ��9���Ǫ?#� {#(&���������6{^u�$(�)�����(������ B�0H��˥�LҤ��;s�` RDL�RG�@���d@�'OP��0��BL.O|0��fDk�'���`�!U���%I��Y�O?*�B�E��s�)���'{'D]P�O�y�� ���;��S�~�k�J!@T�<�I<.E� g84�  b�%
�#���'>- X?���+_�v�x)'�ԵIҞ���[u�<!�M7'�થk�0z6�� �'�pY3��.X�b=۷ �)Ԝ�(��tO��̻y���@lS�2
����T�H����� :e�U27F�٢'�8��I�doI ��AU<Y���3.�O��*a�xbgx�'����עy&D��M� �^ H>��A�!�X���5'd�'��m�Xi�E��ĀN�X;�%	�J?g:�=�C����=�O��G@	n����M��gGn ��n�Cs��&KȀ[���Y&��39媝0$7����gEh�>���@�:L�q"�a:|�xT�'�b HUhXje�͵JM�3GI�2���EF@&Q[�X��$�q�1+1�M]lLB5%�4�Ol�ba":$)���9F�@�#����HX� �'#�]�QH*z"����19D䐤B�n�R�rdF9-N����ďJ-j��&
%O�4��l�6����R4#RR]
��]
n'>4!1^�LYE���u.���P��N�q�=�@�I�"��OJ���v�P�:C�M7!s x�Ǆ�8��">��n�+Qb,�|ZF�_`|a@�R�/�$�3!�`���E�@��,]�<��JV�^^btqP�O�ـM��������c�b�$	��-x�@c��s�4I�,K�qO��$ּ�1C͕O|�9�0i�7D�#Q�A���q�`X38�di#��γm��0�Oݟ0������ ΋7���0уP�|F��h$��bG�E���i���~�!&Ӹ-d8"H�/�݃�a�>�}����
τ�4 �H���I'rm���
p��А"��<n{T���q��P�0�b�?>~8#�@6v��@���(S^�;�uG��5p����r�L��K�=�:�Kf�<Z7#>q��*=|�|R1 ́0���A/)$t8���[��,��v������]��-R��5��Aw(�/+!�D��h{n��H+� 'E;+`��)�M��LB�dx��|w��9-o���-�75�%�E��#�.u�1�X��QSF� ^h�����%4���A�I���<ц#��l��8��֥tĬ�+�w�;gXܫUF�|Ju�G��H�6=��&�Xo�yہ�T�}Fi2֊�T9"��iG�jhQ�Ɠp�H�"b
�\���y��
M{�AJG��.&�X����̝d���$�ܧt�D�:B*5�)O;�y��� �r"$B�kzUS�L��y҃O2X���Č
_���0+�:7�8H����]D �E^P���ӣρ0^���ud,���C�iI�ӧ':�3t^L����D�'r�$���V2�l	Rs�G /!� 9��>��d��O�,6@l$���͓ �����'�ԠRrP/���J��9F�<�"���&�m��A�D *��	Mr���  �?	ɴ��D�P�5mׁI��p0+D��C��B�ZyY� �.�A;Ӊ$?�&A��_)D	�&Sp+�Q`���!H����J�-�Q�`�L!�� 2l��c�"Y}�!���L=+ˈ01�Ç;�$���O�]IvĀ�����eh�aX;�X}(4�.�n�+!O���J1i6>��#k�(  ��©\3��V�<��>�Tf�cJ50!�H�L���^���;� f}�ɽ�l���/�-l]�ƅ�.��B�	�@��i��S�$���	�b��;�G�E�S�	R��x�֖�hTP�G@�8�|B�I��JgN�m1����݀Y~�����'�g?	��K�0�J����L�I��F��J�<3��:�5�L�'� ��2�T�<�`�1�O<mCr�$��qӰh؁l8�Y �"O���WBОo�-#��C7�Q"O(91�o�� ƞϤac "O|��ׄ!&�H��"�:4��|�r"O&���Ke*H��Bd�\C�"Ob���fA&c2�¤đ2A�����"Ob�0D�@L!��c �k��m�$"O�HxG�0?�}:C��-x~xr5"OF���<R>q"T�G�oU��"O�|YV��$OH�C�K���"O��e��jj6}�%�%i�X	1�"O;DȬTZ�u�a���i�jI��"ODt��$4O��L�p��'5�a`��Gu~T�VN8G��l��'@�T:1m�i�
���>>z���'8e�������F�6a�u�' ����;�$�:cB7,Op���'oB�2ćD7y��	8$��$��9�'���P�j�ex��L�p����'G4eÇ�6)V�p�ǅ"�P!�'��e���Dצ�*��:Mg`A�'�$D8�L2p�
M��B�29հ|��'�J�2f�#w���p �9��l*�'�ȹ�����``��G�4jRt��'4��{��*:��qY�/�4$��'��lK�kM� }aq���v��
�'�.Q��n��X͢ӣE�<�*�2	�'�n�pc֍c�����ʑ�L>Y
�'úqZ�`.xv��CIN�P���	�' �5ƃI2�D2@<YЖ��I:VĹ���9>N��Ņ�6���ȓr�i'�P�:�@ň#�E��X�ȓS�N�aச����@f5er��ȓL�`���cMr@W!1)r\I��O�2���y���U��.1�Ќ�ȓ/�xz�e�^��'O�f����ETe6&��|��xՇ��}�޽�ȓ;�����݌���+�)K"��ȓ4����;I�H6mQ�q詅ȓ|Ɛ����Vn�;W��'NՅȓ"��[�g6d^�S��I�}����(�.�
eb��&>����EA�;��ȓ?/���e�<�����9`	4���/Ҭ�2�T�A�%`�1�ąȓM�ƌ2��w�D}YM�6N@A��lM������>�B���m�$`��W����O��.�0"R�J�u�ܠ��g�,-�c��1�10$��,n�t��p��tx�CO�f��"�֒i�,��ȓK`֍¾nL��L��V@�l��5�n�0�ڈK���|�� �ȓ&�\(;u�אjפ�qC�C�Z9~���j�)��f�3&V$%æ8�Ȅȓ6����I�0n�5��=�6��S�? &%Kp�W7���� ��k��j7"On�U�Ջk,�<0 뚦{d��'"O8xj�F�BZV���jS�Q8|H��"O���@��8��G�<+�x��"O�|2��>F���ǜ$a��"ODA����8SJ��B�Jm��m�S"O�)��;Z��@���("�T8�C"OxxZ"J�G�p�ѥ�#-J$�q"On@�J�8Zt)���iF��sv"O��#�[$Nv�!bb�RN�	@"O�%҄d�w���I��P%sV�J�"O�x����~liR���4iM��-�yb�¥8�X��'��H�t�bF���y�Ӿ_���	E���x�!� ��y�N!6wd1%Gז]�qs�n���y�얼f��A���ȅ|C�e@�Ĩ�y�˯&&A
' -h�0��'��y�I��'MZHФ1y�4��W�$�yrb�\T�v�Y�v�"�(����y2l	y�ڥ*c���R�\ �y⎞I��00k��R� ����Y��ybnM�I�\š�_�D���Q �$��<�c���y�T�O��Y�a�����ՈF�%��� "O��$��A|*�`�GJ�|)���>!�.Ͽ.���ZH>�O��k���$���b�@
�sb��1
���	�'����p�G�dz�8S�g��9� �O���.!���K��D�x��|��ؑ8Q�\j�[$��!S̖0�'�Љxa��Z�bɳJ1VV UD͉Nl����h�?�Hs�>��KQ���M�F��Vg���W���M���Jc�MW���䎼)�p�ם>�Ue�j_���#�A*;����DM}B�F����Gx�@�*?ZL)1S�T�v�ˤ�)?A2Fī �	"�	7}���5"6�L�9��S���;�M�BT�Q�"����x�J�>k^m�b��$��u���
椬�O�ӴeZ��u)'�L)�R�'' �]WR� ѰH�-.f,c��A�C��UT������6p�$I�D`}ut���B;"�is�ϓ�L,٤O@��F�>�s��y�S�1c+�,�6j=�0D
w�x26�E&�
U�V�>	��Ms@�BD͑�^��D��Cq}"�V#n�����g�ɭG��Չ	E~©Q������dD-�h�d͈��imaP%�%jGɧ���R4&vXA:$�A:&H8��-��|�qO����O>�DCV�$���[��$���=$�������Z�t���`b$m[:Fg �`��P!����t��|�ΐ;n�np�D����x�F��K��6�FW���Y\��B�N����r (�Pbl�ɒa�M�����Y	
��"jl����J�*���E �+��в�U?�=P��[5ߌA�V���M�B��<!t/A�U��S��i̔1�ʰ�ᝦ1�>U2��N��D9sL�9�IR�R'�� a0O�~��Γ�F�"q��y���m���c�P5��!3��I��$�f�˞93��O�)��;4�X�'z��H�m����[ Q&� ACWf���!�.�*�O��(��f���2;ғg�mՇ
�ie���Ѫ:�2HϓPy����&I�n���K>����n����)B�b�]�R���ZB���f� jJ�`a&ȱ-.���H�>b��X{b�5M�q�P�ߋl�xٱ OC)�Lb!䃇Uf���N�􉔂���Q-�.?�A8�cD�N%�|��
���Ǡ�6[z��� C#��LIs�j�'k��o@�h��'?�P�OA�h���/�.LN@1c��6_h���ɚ�B�-J@\	*X4Yp���i�
�F�>���i�]�5��:=�a�w&���x�@�^_��Sa�v�D��J��( gǃ:i��L���s��S7~��ԥ
9<y��Z;!�,W$
$E�2�B�E[4<��O��IFzB�0c+`K�� �%JP���y��ֱ� ��т7S$�˓Z� S�.�	�V�p' G	,��	H% :X����F�KF-3����W
����L���OnH�ꘂi�B �a������J:Vѧ�ƬYYd�'I"���ޭ�~ey���$Ei(����I����+�׼ˀc֟S��H۔��VJ~�J��L�'�z��1AF�;��%>�jQc^s����M�'�n���h�6��tS��ٝ8�ܘ[��O��A��	6g��թ�n�x��?A� �Jxf�I�∟Sp��-��XŘ�v-��'���_fơ�'�Ty�;$$ȭ+�JM�(����2f�}^B�Sb:r��\�2Z?�2�|>#>iE,�$a�&q��X�uezy�U��p?iW�@ʖ���Kn~�.��Yז^�^	ϓI�\EH&��>Ut|��?xT���}�� �'�f!��B� ���
.�m�)�L���EΜ#$;��{6iU�fBv�'Ir����r>���$��x����D(H�G%�O��0gH]^�? ��j�
Sn�*t؃����@(�B�,3�$�&�"}�;]l��	89N� �"J�`h����O1Ȣ?1%lЃi�*c?}3�H<� �۵�Ǭh���Bm���#g�q����X Py�d�_׸x+V��}�P�퉗m¾L"c��(���Q�FBl�4�
r��D���N��y"�Ff �$�, "r�����'�� �`h�N�E��K��}IE$I( %PpbҀ���y��lS�kv��6}�	ZQb��d�q��=d��X̑>��|��a1!��Ai �^�H�FH�ȓ�J0��EK o@8]Y3(L�[E
-nډd=�Xi$M�&)i�{ �	a�qa2�T? �e w�\?�=�G��	�:��'��OL�X�'�x�J��a#ǺFנ�"�"O&�Au��j0d�i4��}hH�T����� ����U	�h�v �s���2�����y	�0��"OH\�e�F�*��`Q�]O�4�[V�Ą[�b��R�|B�ȱ)��@p~�H�b%X�}�S�8D�l�-A,4K��W�f�"�Qét����C�EI�|��ρ��1sK��F��P3DB�y2�qO<��k?iԨ	�#��y"D�8 ���3���db�i 㓡�y���k�uYgN�;
SƝ*���yR�&2g��� J\
�%	�eԥ�y�O���ibc(AI� �������y�i�E�~}voM1@f8A��KF��(J��W��0?�6&�;j�0�l�1�d�U�R��d.7y�ȳ	�<�ōV��b��A�T���)t�F`�<�hC_l���X�O((���h\?�B�D8T�Ptj!IM�F5��B���ۆ9Ҏ�ȳ��3J=+*I�Ux!�$�? ��S� >�|��@
�*�ٺc�������>L��� Fx�e;_x���_I�tMsu)X8��>yU�ع _x����I�U��u ����Ba�d�K1(�|8%�߅Sj\���X,�l̢��˼�x�ڕ���OJ	��uk�6i���ЌZ��h��ӟV,J�
��g��#F�P'%�ĕ��"O���,�Eլ�H�'P'M�iJ��'θ �MK�a}i�,��a�����33�vE��[{j�yf��/*?\��8��k�o-L�i߫4��I�A۸2����Đ�V��b�	v�d��i��e�&�,o���G�x=b��D{7z��vO�p�>03��]C�$)�FN=�L�"��1U�����(�O���@h��f_D1��fǾoh�z��	*r9 8��XS�"��q�����'}�t�`Ӎ#~�����+LpF��ȓ.2:E��)��B����̃8@.��	$.�ޥ��͌0�� ��d�+50MF�IƮY�>�)v\)�I���C1?!���P�{�%�% +v0C�-7�>X٠%P�eZPT"��G2f�P�?#<�+�j��ȣu�����~�'�,*��C�.G&����d��A�0D�vp�K�RKҜ���YW����k�-<� �	���1r�������7�%f.��L	�e��J�K�`D�A����<D�X�c!W4����M��@v&�O���Q��~B'��2�(��=��b�	<�F����]=g��D�'���B̻b��$�D���P�iO32�"Y����&!��G�8r��aa�'��ŸC��#u�qO`ԉ7,Q�r9�̙����;������-��}1wN�8�!�ۢX�V��E��"E�V��ӻ_���i�;[6�v�ܣ|�'��0)���~��PA��Y�,��'Ze0��L9E�#F�$ 1~��e�@q֤� ?�0>1���^2 ��"B�$�"�]P��l���2�A74O��b��N�ε��*�p�C�*O���qo4�h�ԏ��ipX=ʉ{b�5=�ո�n�L�O��eє��7~R�[ě81�Tt!�'s�qا��`�d J�b4�H9�g��xdiN���<q�H��X�"I3�ه]H��(�S�<q�	18b}h� ��le�t�T�c�5	fǀ-�l;�S���6D�r4vت��0:p���Zq�u2GNr?q�JE�F���+7�@'$�-��$��S�? ����3/T����E�5DH|��#�$	uy `1���Ű$�@U"�&~�p9�!K�.�!���|�Z]���3�I2�$[�!�D�+"�v*��I�w	'�!�$<�.��ō٦{�nر���c�!�d� [�!pR�߂Ri������"�!�ā#6y����/j�QSq��!�df�r͒�0aP�e1�R?!��[Ů��#BJ8%���a��y!�H�P��k���&�PW ��U!�dȻ]NE�A.Uj|�$�d�o!��8m� �b��+k&�Y�i�'!��Ѕ>�tbg^�6����t�Q(!�DX?\���k����?����vC�-4!��.��]�g����!8�M�R'!�D�5Nz�R6/��6���!nK�I2!�D�d�9y��#DɊ��nE�C;!��O��)�c�C�
����RG!�d�d9� I��P�#��qX���1X#!���
94�4(��LEf�I��߫`!���O���ؒ���p�܃E��F�!���OT�]R���3�ah���\y!��3��!X�
�"�P9�1�S�E�!�:P/t58-׀�0���
9�!�䋠x��1�&��*�bJ�aλ�!�D ��{g!I��:C�툧Kq!�d"Nι�5�FM�*��DJN�Q�!�Ć7K4����1x�p��X�n�!�$�^v�:�R�T�� ���1�!��7�4p�I�LZ�=�ǂX3w�!���L�����(\1�E!�ܞE!�dŧV�LY�Պ��|��Wo�*W�!��z�l��`)�J����B�[�!�D�0%�v��e�L����aRgI��!�9S]B� ƞ�ݲ,�%?*�!�D��r��R'�"\�uℜ$!�d��X@���W�Ղ80�tq ���2!��	��08�W�z���i��OP!�QX�`qҗ���X��q(�iP�]!�D��C���X�n�����
�2!�$W��t��2�Z5���c�(�L4lI��,�a~r�� s'шc���Ɖ��y���lm�"r$��0�������yB�6*��;�-Z����%�yB���}F`�ڒ�V��������y.���5�SJ�vX�G�G�y�F��h�H��P�&vQf��&�J-�y�S����ɝ�X�F�1Uk���yrLē��8���%D$����E��y�	R'6�8aZR�'�$��G���y2!�!	�p�-�&�K��C �yR�Y$;(Р�	ŠT�
����y2��W�V�s�*P:L�D�`��H��y�D۬�<���I�z���������ybʌ-mmT%PL�m�����/����=ٖ�HN}r�6���$�K<���AVR&c�ʩ��A\མ�o�O0+Dn]˨��Eʷg�<Xǰū��G�m�̨�G+$|zD̋e,<[z����̺z�����+���6ő+6d�x�R�?ߘű���/hR��rc�I"����OV�a���I!n�|kԣ�� �t8uE[�m���Ƌ�F<�n�0|Z)��p�`Ȣ'��2�p�
�#e��\b�iX����B��\Ep���i����ɅRɪ��h5ZY8�H�P�đ�j��$��?U"2MА{�����+ȠYN��w���؛E�L<^@�$��}��+qu�&��1G0諴�T��h�G' .hɧ蟾<��g��l�E��n��#���cϋ�{$�O��k �π UCs���4��p	'CV0_<�MAt�1�d�_=�IId�O 8�3 �g&�ak���T�(�'<X$Ia`C�Ć���7t-�9��'���@EƖ7}�%HC@�Z�\�'�P c!3:�T�b*ٳT�>u)�'�aCFl�CvК��G!T���H�'�W��Uv��$,��-�#�N�yG4 #�0{ g�)Y��*d �0�yb�	u�&M�FJN�'�"�I%��y�`ƴY"ǈ6w���	�	��y2*ʭ(6�q��ߝsX�
H��yBjۖv�2��2!O�Z-��H��y�/F#(HL�b�A%FƐe�Ӈ�7�y�c	m�x�j2A�9�mj#�D#�y"��IƂ�h���C���֥��yRW�O�
�1Aɓ�A*����?�Py��߂��u���CJ_f�BV�d�<)��_q��� N2���"�u�<�#�N8 Uz��`O����r�<�"�4���š�d����sG�l�<a�a��~/�%JP	��3�����@�<�bB�.n�)��GC4j|<ɖ��v�<!����@0W
ճ8�,d�.IX�<	��f�\��4��-7��H�J�l�<q2K�3�&D9�(c4�@+�^�<�r�Ź�>8��E�XR0!�%�\�<!�g�iq0�0�64I:�.�B�<��Si� ��k�:G��u��D�<���R���HA⭂��hiʆ�BA�<Yfj@���Qi�[�0��L�h�<!�ַ�� Bӟ;;�Y�i�<���T�G$`���L^�D�>����@�<��^"I�,���ٓ�0�"�ɖx�<� 
J%>R�0���鶕���Y�<12�Y2R^T���֧0��@G�[�<�S�òVd���/z��EiA��<�'���^z���(\R�<�7� br|��C3� �qWOMP�<�b��X�Ҕ0�*YU&�Ib�r�<���2
T}�`K����0@�e�<]
�;O�� �2/��p�	�'�x1V.��;���x�.1/|���' ����(�>�5ۗ�猘��'(��HR�O'm/�|�p���i����'v��X7a�#�T�a�we ���'MT��?*w�%C��t�0���'!�m�'+�.l�rY8Ã@�u{����'��P���ڧ<�r4�-� ��X�'ژ	"�e�{�F��%  �'�H��f��"chR�`��S� z��'��x������-k鈂1�%f"O�غW�;����(аcj�@	'"O2��G�Ě$0i�Z�7&���"O� ����r`�E�rrƜ�B"OzTcWfގ��8S�l�I}�Y�%"Oމ��g�E]�� ��1do�	��"O
����ϕ&��Jt$זb
��"O¡kV
�]t ���c�0���ɥ"Oh�&�Z#3~� �B�(?�\��"Ot���]\�p����	@%"Ol}�w��{�r�Cg�D�� 蹖"O��C2:\yX�D�m�h� 5"O<�����.D5C�C�$Q}�5P�"O��&�S�pQL��ec�eP!R�"O� ̽�GHX��y�!X+�� �P"O@ '��H��*Q-�� �"O���+Y% ��Y�O�)<�ܱc"Or�҇,!G#���E��F�I "O��["JMe骙z��
Z���v"O��"��sn6��ŧ�8ui %z�"O�-��	'�B�kR(ͶN�J`�"O�u@&+�":�N��%�����"OR�{���1	��L��B�H�ZU"Oz��Ԃ[�m|Q�!�T�R"OD���&�s�d$���p��"O��0p、�V���ȟ{�Q�A"O�8ګ}��AˑƜ=���#v"O��sc�fZU�@��<&�4�C"O�zmc1*��]N�@�A*Q�!��j�f��GB;[��A�
*^�!��[^�]I�B4��Ɠ1?z!�!"U�ypGm�-_ �[s��%S!���2Z��Cj�T�Re�����]T!��J#-c���j��F��Ųe�D)tO!���,� B�9&Mv��5�V�X�!�$�,m��4�p�K�]� �T�!򄈌ה�yrF��Z+[���6�!�䜊މ Q�S2�
�Y�.]�"!�D	I�Hi�dQ�^ņ� ��Y>0!����pe���L���g���M!�L�2��9#&� - ����w�̏B�!�D�]��lS�����"�$R�P�!��%g�0���
�ly�LjV�Y�i�!�dU>m�"��׌\�̱V��#�!�Ԋk�����O�p���҆�~�!�Ć?��e�d�^΀}��ea�!��؊������/d�D`��%�,!�!��m\1�C�Rx��!�,�!�	�`����h��`*�z�P�(�!���2�X��fM�9��*'��O�!�
�!��� �4�X��v!�	U�J����I�0����b!�M�dp �c�3���T�0xo!�59����	�J��S&d�=!��7u˘���G:2jСJ3)�[�!�C"(���p���
\��pR(ɐ�!��+6P�g��c��=I��P�c5!�$ә%�<�JV��A���åA��!�DK�(�H��%��Z���I6n>l�!�$�'YcIa�:/_���mV�[>!�Կ=�j���[�uU��q�L�1l;!�Mi�������2�ȣ%+��T!�8H���I5��	ij��Hc	S!MB!�V©۰(ڃLX��cd.	�!��ڹD�1J3H,u쉩 �D?/M!�$20P��+�%PT�R2RQ!��!I��E�u ��hI9��J���Pybm�/��]Â@K}�����	��yc՛)��Q�T�K<0S���AE���yb�0]��X���S2:i.@��(�.�yr�ӽNxI�qIͺ0�R�1�⚝�y�cV�_� ��c�#s�u{E���y2&ąT2��q��(;�d�e��y��m��	*��T��  �O��yL?C3LTC4�����������y�'� ���scC8yk�[r�R��y��M�I��	a�R��������y�c7<Lr����A]Z9��^�y
� H=C���0s"�3G��L0�ى�"OͰâǹS��D��[�2-D���"Od����F<����3|ڤ�A"O��ɦ)	����IM93�f��"O0tp� `h�8�(�3��,��"O�����QV2�`#��6|��"Op�XnK�,⹉#����$0t"O`��$mR�C�8A�v!+lJ��b�"O �S䀅�n4�-�-.T��"O���M!:"޴���G%��"O$4����<�8��0b�'� ��"Or0*cmV�4� }��j?RDv�
"O�ق���8=���Å";&�s"O�	����X�A���E.�:a"O�P;��G�>Ԡ��B�P�;�X��"O��A�֠>M��s�L�r�옗"O�!*U�D3�d��^ Z�&"Ol���IMC�$`���0����"O�*�O̷��eiP��!O[���"OH@ɦ��=P�c��\�ZWt(��"O��ˇ��@�Ⱥ�H�	)>�"O6���lmz�E��Ȍ!2@���"O"�Qcϕ=8w) jۉGQ�p3"O� 84
��L�ȕ`�'TR�eY�"O8,x�a�l��hq�=5;n��"O�:��Q6L�lb��ݭ*�M0�"O��X��#����r��t��D��"O�MSA�E"H=�R��Jx~�1""O�����Qd��#���eЉ��"O�X2�����8P#�.;6q��"O���:3�*챔AJ�n �S�"O�Ca�V:1
�` =�,���"O��6JO�*��`�`B��-�0"O��dł��!Q�/�7}ܴ �"O���H�o6zh�6oK7_��Ȁ"O*��e�D)9x�`p�n:7U�}��"O�l��	�Ug���6��.-�;�"O�8�\g[H��#��9n�%"O���d���S"U?i�&Ms���y�V�lX���\�r��`,К�yR�;K��@ٶi2�\!�`���yB�ȶQ�F�W!�!U��X L�+�yR���h	B�&<J(�(
��/�yr�R6�
�8͉)B�t]I���y"�Z�(�XZ%���9�\����y��	3��Ͱ�*X&�:U���޲�yRJ̬k^\\�S�3~8�Y{�����y�-�`���P��C�z��A5���y2�F�@��-��9�xUo��y⇗�=1���T(XT�������y��>|t#�FƇsl��kN �y���7y�V�9C=v�S�V��yr�ƈf��x@�h�D�:d�.�yB*��"MB�J�gĎfY� #T����y�U�}�0̆�k�1��Ӎ�yb��L����M�e�>��r���yr_^�MIs�X.t2Ԙǉ�)�yroG�*Qq��Ѥ$�M{p���ydEn먹�Z/1d�!�4�ۺ�yBD�46���t��N�Q�	�'����d
[�z��5�� 2���'�:�f�߇u݄�!��xF�Q��'��	�%8v���ԩN�mMA�
�''�`���<2o��b���)\9Tu�
��� 0@�D��.t��"h���J��5"OD3&X�,
����ϗ�x���"Of�0�G��"�$��KP8#e��*%"O�A{AB�d��P;$,N�"tZ��c"OP�g�Z_�HK��D��"O�l�A��c��$`�6�&E*G"O �C�   ��   ;  �  �  �#  d,  �6  �D  �R  �_  Mj  �q  �|  �  /�  g�  ��  �  3�  v�  ��  �  R�  ��  ��  $�  ~�  ��  W�  ��  ��  (�  g�  � �	 . � � ># �) 0 ]6 �@ �H �N (U k[ bb �h �n 1u �{  `� u�	����ZvIC�'ln\�0"Jz+��D��}�2TP���	#Ĵ	G���?Y����y��2+�<����3:tE�u���WN ����3z�Z��PI��Cb��Q2���YYV�� ����WK�X 횕2���9�QPr�WK-p�ݑ�$ }�����K5Y7 l�;h2N��'�?�⅃*R�6�X��:!'BL��>+��K�h��e�r��ObH�FKp����[�^���'2��'=r�;;�.Ժ�fQ.��m��ϐ~"�'C7�P������:��X�I+D����۟(����S�D�r��@W�� Ǽ4�I��(� �X	�fԟD� ��3�^�韘扟@���ہ��Q��x0#Ǻ8����F�: L!�'PB�a���o��p&#�",��y���	��q
����ͼ�էu׾���]��� �ó>a�c��J����q�S�V-����!,���Q���?���?����?I����'�n)�p]�n�@���n������'}�7�Rꦑy޴OR�6�'���Z֍rӀ!oZ�M��vBr�/��w J�a�'�P�4�'!��~���@�r_�2㢘�t�\`r2D	$z�ደ���(���5))�x@�D�9h2b-2��@�?�F!�Ri�3�.��]Dh$�4��%&�+eM�!������f�v�K4eH��E{��Fi�9��B-1��l�c�] LJh�2�)%e����/UZ�Y�D׋X.�� �I�B��YI�dͲC�DٽK�|0s���1�b�9��B�[�N$�#�9`T��V��!C�M�G�?!�ؠZW�+I�����H$_�a`lBu�: ��B	��*���D�G���9 h��kLr�0Bj�r0r����Z�⃋B����;Ve�k��d��%�>m�-�"�� V �����{|���&� Մ�0�#3l�L����9w���&M�c1�!�s�\�L38m���?�{�'��`�r�c�m�ןj@Mɲ���$��ju��v�Z˓�6e���u�dɎg���%�;�	Dk�l��a��q�a����N�axRF�E�t)���|�µY�9D��N��ROƂ�0<���]�����P~F,-Z M��זi���)���?����?9���I���BQl�$R�.���K�p�qOL0Gz��"��� �=B��UIA䛌o�=#���l>��?�ɜtw������ ���%c�j�cq"�T|V�Aよ�2��'�Dmq�4��x��U&��庰c�
*��l�!c�yR�H�{�2(�҇��ue\������ē�hO���]`:NU�8Ap�O�<����"O�ш��Vǘ���)�����剸����d�'�lɓ��ա}zN=�b�M�VӤ�S��ܔVT���<���M�O�^��'Ő�c�$��1o	ZꐌB�i�/��a��'�F��S��X0��8RjŵJ<��)
�'�J���(�r(�T���A :���ӈ}�'v�Yਫ਼8m���9�	G`htj	�'��q�b��46d�<K0�ܡB��-� KZs}�J?�.gqO���J�i7*0k� �Yw���&�'�(�k�L���';p�@����'��i�FԉM�b�F`�>S�xP�D"O����@���(�լ4�O>�(� \#zHvT��A�
����"�W�<���޺%��E92�ћ�f�4�p=����tD.d�LP� ��=[��bqO���<��FQͦ��&��x*���,�ҕ�C�kc���
�<)�	�X�T�O���MD7�N��t��a��EGl�Hg)�:gԠ���'8쑫!,ª|��'_������ R��٣	O	:��[�L�����ǟ@���P���$��8��i��&.�x���\jy��'T�OQ>!�j�=�=���Z2R��� �HO���;�,Wb�:Pj���B���⟼�=Q0ʎm�1�H���,qމ{�oP�@W���������݊�1�d��I��!c�'���K�%3ZyH�	ۈ��5��'�(�4��D���i'������I<I����ڱo�
��B�$��ݸ%ϓ�T !�䊈��`*`\�(�D�&��Q��*�Op�Fy�����h��ft�s�b�7Le}kH>�F ٿ-u�$�|ΓS�,H[` Ϙl��!�@S>q*������<	2M�OҜ0m.<O�}��Ԗ>�pd�&��3u�*�X��ĕ�B����$��s1�hb�e�&�Jeⷫ޷/P�����N�O�b>���O��d��0���
vJ��_i8�B6��iB
C䉏T�����ʜ:�ȵ��.���!6OP1��4�8���<a��1h$T�
 ܁"�XYkH2ޤ{f	�0��'"�A���
���	 �hu�t����8�j�n�s0��(�h���H�8�Qj�EtF��sÌ:[�hB�	J��(A��X��L`��,@jU`��O�!��Ɇ|vę���	=���P�0^Q���ğr�34��Ku�:�M�0*W9��L%��H�,W�I7<Q|�A�#֟p���W~��Sт�<|3�,K��ި"��	��(J!رVZ��IП�C���'`��3?�� n� ��ãQ�����
^��'O�)CX%b���g鐠�yb96�H��F�J>f�S+��0<�g�O�,����$� Kl}�@�)\� ��2���'"���9�ja��^ՖQ�&�K?��D�BC�	�����&kfr��C$�cf�a��Q�LJpȀ�Æӟ�'� 	Zq#R1L��'哖&�F��=�0� 
H�?V��A�T�6��@��П亁�6tҚ�C#��Y~�'V�@����Pjt$
�a��A/Ӟw�(a��h~�н���Z�e��0|�
*��xb�O�v��͋[~��� �?Q#�i0�6M�OH"|���O�Q:��H:d����C]�I��(��	�j�8a���s�M�#ϔ/��<�G:OƜR�	�iؐ�q�@ep��1AG�f4��V�ܟ���͟�h�@�}ބ����D��ȟ0;0A�(`�ء�)`�pi��	�6�E�4?ٲ�.�0=�5��
UU�\�S�R�0��K�e( F�(כfo��M�������y"�ƅ.�� 駯K�R��X�(ִ�?��_�DJ"/�Oc>���O
��H���¤��N\ic�/��r�
��:���@�ڱ+�n=Y�:���G�F;�(�v=O8���.����$��I�?�'t�պ���g�� � )�Y&�5Rp��nT�b�$H�>VLy�$�>���*e=t��&y��	
kH��Ձ����>iWg �֕�bB�RƌjDm��(9��@s(����>Qc�
�xw
�0���:;Lf�z��٠@[�4�Iן<�I��'K����;����$bŝ^hр��U���zܓ@�
S�(��1���v�O�$y�p&�D@Q%ߟ`�=ASH�-C��Ӳ|�h��v����kƄ-�	�֒���"扳��>rńS�-]u�Ǫ�T�z%��>D�l�S]��e{`Ɲ�PonM�F�<,O�<�C�9}0�hffZ��Z`ҥ��q�<U�N�b�be Ҥ6v:F��2��jܓ
O���'P�<�0G�*}Q�jX_;h)�B�3�#���r��D�=Z��)N-/�H�a ^�G��8P��զ>��'�lA��CԎ�p<u�D-TQ���%�j���La�<�R� �7
���Ǟ|��I�EJ^��I���Ot����)r���`�b��0+�'JF5+7dZ��H]`��^�~�3��d�x}��)ʓZj�Q�ځ5��B���(�\��W�:nVb�H�6�.§�>Qps��7d�j��VJ��H f��v4�I������lV=U&���6�G�kO����%:N)�E�g螅�0hA�0���>	דL��<ȖE�Pr���E��5N+|M�ȓ"�n� EN�oe�<Jv��;���"���W���q�{��2v�����N4C�$�R ���?��O�p��<)���p,�y�<a��(1������+4C��1)�yB��`�̌����u�&dZ���3��x�X�N��x�)G74Ǧ%J�E	�ThB�I�!�N��ċ5��[b�
,�����P��fL��呫1�n�"vM�	A;*��=y��	-��S�'kF���$Ҭu�� �(J	�Fl�/O�����41O�qs�)�>h*� �>��pR2�J<X�!�$��v6�Se)��M+���T��ay�I.{b.{��&�f���]P�C�ɬ{vE�f��+Z�d)�W��V������?���(����æ�A��$�G*��N�Q�X�WN���'r�)�O���m�(9m���ܶA8�K>�cc˻׺��㉨~�� ���`��@a��l~�B��0AL¡�ɒ6ΤȓaΘ�|��O\�=�~��lϖ�~�����;�r���WO�<i"�Ԗ>���tJF'Z�8��0Dr�'^H�f�Q��B�H�> D+c�>�E�>gT$-{�D�{�>��a�]�1��� Z$Ԙ��ۨf]n���,�؁QmDT�x(�" s��Q��<D�B�L�aGN���)�P����H;�	\��<2��	u��,�`��-̀��+6D���JI<i�$��l�,.H�� ��ɱ�HOf��=�!=_�"��/��Y3\���s���b��x�V��c���l�.;�x�pD�.#5Ĭ��m�<� Z�3O�N�0ԃ2G�_u��rO��s��[B1�H����I�*��a�t�<�T"F�K<5jÍ�#[pt��1�e�����{2nK'j@uВ��8����@���'؜#=i#�L���M*(�n<8D��q4p:i	9Wg�I-gר���#!扃4���>i����\RL!�JI�j����=D��	W�؁M�Q�+��b�a��;,O,�<W�5཈sϗ&8
�`3eI�<-��r򅚷}�.���KG����=�6�):�攗'ubň4��2/�%��$Ds��<G&V(X�1O4Ej�ן�1��	�����ZG�D���|B	�'G���	Ǔ-�P����?�@�;Ǧސo�B5��bb�\[�$�@{��;��dR�$��D{���%J.S��`@���vx
��V��yB`X-Y�f�H��)�Б��/�(O8T�'���<�[�o��!�"���=��MRGC��\�0i!�ɩ#b"|���L��Č��e��9ѰmX��\�lS���D@	](<qG�nF�ͪ�ML�BeR�9V(�]�<)& M��H�����_�9 ��_[��p=qa�e������S3p��s)DV�<t'�{V��<^I��6��A������ډ{B'�����XՊT|�=+F�V�?�$!Z%*R�8�<�q��*de�<�@��O~$(ؓ��M`���G���y§C�Fq(� ��{�R� T�A���x«Q(a~nl��aP�lr,�_�eZ]��'\dp��eA�K�(E�����=�{"(X6tƠ�����Jn��G���'a"=��O��5��Wi�ȸ��rD�L
�1�剗|��ɹ1�I�Yhb?�a�#~�	�e׹[��Ӑ"O�t�f��)d�V�C$۹x�i��'Q����a�Ld
m�>��)��(D�l)FH�_^PI�Q�W�#}hh`Wi'�HO�Ӆhrx���)�JO<�@�%\��剋O߆�y��׀��t-(o5�b��K&5<H�KpI����-�*eH@nAc8���U�X�[��؉�H)F�� �3D����"PS�!@���!?�d��N1�<�S�'x�`4���<� ���{P�d��l�*P���a��I�Պ��5�pXDyRf�>� �	�k�C�	�5\�<��;�8����I�`c����F,�'3Tjih%��n���A p��(�a�+�4���(c,�#�`��6t�r��Ämf���)7��8�`U�y4�s���W%� �>��0�6��"O�&6*��WJRr0��P��b�Q,]���@��ZK�D����>�3�ɳҸ'��8��^y>w�ك�B?a����/`��3��>Du��sU�d+%`��(G�R>z���HT ��;P�C�	Jz�,�E��� pA܊C�	4;�vI	��#l/�1q���^l�	��'�&)�	�Vs�TQ��*[i����~�qO��C4�/D���8��[���5#���\�'��) c�>�G��8	q�����P+>��R�(�<sfC,���<��	�'S����%	7m<��I�&ݗ#0 ���C8�1���搀�p# +�˓�(O�ء��*9D�	ANV�#8f��"O�ѣ��~��pPw���,3�V�ĞP���ɀE�"$�	�eX�aHD$R( ߸L;��Z;,�u�<9'�i��G�[�*(��g��2
����d�	�'ݬ����:O���H	e� �quFĿ
�A�0"OD��O� v��,Z��_=��bǕxr�)�ӑ�pt�ѐ3�X�JC#�ѡ��Y@@��S��!|x1K�dW�	Q��`�O �FyR	�������Ì#��
! ۚ�r-�g`�a�>�h!E���_	���KM��6���cǭBNаfdϽ�Px⢚�:`�`z���a3@��y
� ������6b�����ɖ �*�����2\O�H�p�M30�u�S^\�<��"O ��g #�=�$��J�B�QD���{�'O:�����0^����A�F�D��%�O ����Cp1OT@���<H�1O��ȕ.�	~3��-~���4-0D�d;`lIC�ڷ��0m�8,9��.$��["�;_)���B<E`XyB �ڑ�y�Fċ4�8���X>���xg���p=�p�D��6-��c*�#+q�X`GdW�R�qO&�EzbH�."f��ɮ
1z�:��N�$A��tl�:#Ô˓W�H2s�Lc̓���}*`��!
�����/ޙgY<Ѱq�Bn�<���7�T(��I0��� @GhX�LFy+98��& �	V�`�����y"��>�Ĝ�BH�C��]{�JI�'� #=�O�^x`6��g$�"CS#Y����Ox�'�Ly��!�	$^�^�'#&����ym]�H�[�^�O.��#G?��x"D�Q��r�˧xQ�(Ӷ�^�y�	�!1`�ԑ���^=H<R�	H��ē�hO��"������e��JA"0c��Q�"O���gK�"q��)P�ތ;E���ɋ��d@�'@>P����x���qv�KN�<����7��<)Po�O&�ar�µL�a1�	�c����¢H�*�;�'�
t�V���;��0A��pJ�'F�D�gb^<P*�l��L�( �}��'l��*�K�.���1 �+@� q0�'�xq�nB�	T� @��5<햸�!�Q}I9�pqO.��2�E�)�Ay0 ��|��٘�'���g�+��'�4��g-��֘'36�F-W�Sؼh���X!�(��P"O��ӓ�\��4��#H��rO��Ğ�z(+��Rx<�\�C�{�<�")\+c����M�P�gG~���I�{��	�:0�5*�灧�e��B��'�b"=�*�2��E�S���ɂ^#���7�Ȭ��*"F�X�>�s���>- �+_���ޜB�*�z(5D�@2t�M��l�Q��ݰ1zf�%,O��<��������9t�C�%�}�<�Uj�i��1�R+Y�vD�ǘsܓX]���'Pː ej�Hr�=�G�O �p-��:ʓ$�R����D�g����,MՎP�Y���4��8��'�T\3jհ�p<���<k �\Jtn�!0�0Z���I�<���r�@���~f�h� �G�	@���O6^�����7f@K��;sͰl��'�b\�����~h�șn��?��U����Z}rM-�8qH��^�lH1��	��d��o�8K��b�0`�c$�'dP�1�@�ՙG�����Âp��x�I�<Z �7�0�!0��-�p	� �.L�l���Jb�}��[!�p<��j��q�D�>�ד*3���\ r�;�Gֻ*,��@M
�p���&Lf4���3HP~� ��>�F鉙��'�rT�� ��Yq��I�d{�k��Ɓc�H^̓g�$�ar`�j̓zPHS�W!M�, f8-�n�A�''е�4A��j��M�b��:�v�b�'i*a����1s�,��`5��Z��<D�ܐH��kk1�����Lء���=\O��=����P�nD��A\�r��1��Ivܓ� 0cX��~RA�.	b�}���@�eʼ� J���ۂ!xBL���d�}*q���[r	��tu9@��b���"O��Q����>�FGӂrT[s�'�Q��A���x��!ǘ�(�Y7 &D��Є�+m�J���F^�
�Y�o$��HO�Ӡn�Z����V�.!ʄj�I�F�0��!ʓ	T�I	����)��)R$'U��W�|c� V���';���P�	�p<񴌝5FH�닟W��k���y�<�(������'LT�����~�{���π ĉ:qf�10�>M+2f�1BΥ��"O^$���rU@��@0���剏��D@E�'��]r���8�d0;���^��g�ܜxr �<٥�T}�O�n���@��J��ġ��ܞkR�)0�
�Y  ��ēH�q����f(�h�oU�:��<�ȓ{)x(�g-[���t�7aLa_���>�דkxq� �t�芑A�BД��; ֹ#��[{9l=�e�|�6(�#͹>��I�۸'���P�LߎOhh���¨!�(����)v6��kYy̓|$�5����}�e��ȁWi�Hf�EMK�����'�(L �^�5�(c�l�0n��
�'��k��}����IQ�TIؙ�Sk9D����U9W�H����ΙX�j;\O�5�=�sj�.��Ap$H=Ĝ%�Zqܓj瑞`e㛣�~@�'��$�í ;L\�e����d?M�������<R�q�й���� V�%H#��+(�ZQ:�"O�᱄@ͶEmĤY1�Y6�4����'�Q��r�'�V�`qS�,S�kI:ɐ3-D���4LG>6��œVc�6
�Z݊��%�	y���iQ">
@����&7;Ŕ3B!B�����ĕ�w����<� ��C
a��1\*֕��惋;�*��Cg�C�I&���� O,�xf�U/	����$��|	"�C"O�Mi!cW�kX��B$ʐP`�c�xB�)��n츔���Ot�t�(��\n��C�F��P���
=8F|c�eRv�<y�X�4���$��s<�D8@m�:<h}��	��36̑;��'��b��IM�+�xAtEF"0	> $cԄy����pB^�%\�𤒀G|�����K��lY�jC��!�DD�#I��Q�E�-&r�!׈
�n�ON���زD<B�!����"�:�@C�N�!�D\����\(:�& �fb�	R���*�OP�Ez�3��ENA�f�ϡX��,�c��B�RE�����O�3fCA�<��1�]�Bצ���'�f�[��m�g��y7������ 0Rp�<��'��b�� ࡏ�]_�mY1��O�$j�	P�*�;�c�_#����m��C�� *"mV�H'��c�H(G�b��O\�$O�;�F�	���!d,B����'aR�'1����%ꗪ6)�� u�֥5¤qP�]���I}�x0"�Ц:H2����#@t5ˁ�>}B�?�S�TD�-�~�1w�hx1B䜎k��p�fL���xs�Ƃڋ-�%?�����?�I�[�^5Y�㑍gݴ��c��1���IRI`�a0��+qj��2«�s��퀘Z�	I?�:��B rH�D�H�1c<�y�YGJ�}�Rl�b	7HF5G�t셲���d�J\ m�F�y�Q�?1��������l��jZ�!��*�	k8!3K0D��1 X�P�h�'�'w���c�;�y2�� �O���l�@�58yT���ɚ"����O0�dՓM��8A69�P��Ov�dB�{���G�c�r��EkC/t覡��hМKbF�2�O���T�*�z!�?#<)���)`Fl� ԋ4f��b�e�e
�	�1Ռ@ ���>�z�g�'I����CN�"!��h@.Ć* �Q�OLlC��'��	�<!D�+q뾽��&�-_r�rG�^@(<q��թc�ȅ�G�~�RȖ)
����>`y���Hԟ��'��YX��}�����jE�gLn�A��n�A���'���'�b@�'!��|HR�'
�	
T��P�7)�0THpAk��L�hL��i�|�~�+��Zl؞,`�FŌ؊�B|�60rTg��2��h���(a���ۓn4���I%�	dɊ8-@����H�^!`��I\�'w�0;0��b����Q%M�|d�d��H!OdaFy�@5�����1� �#����$Ѥ���$-�I+y�.��O?��0��F���FH2	��R&��O�iK۴(��c��
�)�']��p�CM7iB��;q#�7Ӟ`��'�j���lƁw�
}ijC�'��Xӏ��2�'��0Ԥ�+"�yy׉��$mP|�ȓk���B��\	B�ɋ/�HU�O0�Fzʟv��u�L(f�Q�=��D��G��9�=q�d�=u1O��J��~�4!���*�E�˓{+�b�<�(P��x��[o��H�q�
tDv�PF`�plx��'D�`2K��y��,�,�s�>����3� ^D[d-;����W�
{F`0�"O�}2� O�eƖ��TI��o�AX#���w}��2ғO�c�%ƹH�*��U�Y��P��*Ą)�1O�P��;�S�==x�aoE�bq*�#�.��`�̬��H�0�<ȅ�q\�����k|dibҥ��Ӷ̅�I���0��Z'�4�(M�]i&0'� ��I�L4�r4$ :=�����~.�C�Iny���$CI�:�x�Lټ"ވ��O��EzR`.ʓ�a�f=]���!΍c������)��c��	��ǩ(1Lc�k@+ҩZ��h��-[�y�<pʢ-�y��`�ȓNUl�2�&�+#��QF)��Ll����Z?���
j�1�vNM�a��Y����C�<���O�`ʺ�T�?e�eà&�8��2��ċ&x�v�+��H�=� �g����Y�1O5��m��$�O��ӒPI�H"�h^�h3�M��#����d҆B.�9����O��$��B�C��u�>��8L)�B"�֮uA%�_�GZ��F|"�M2\(�	p��l�'D�L�c�<�.)Y�NF�F|�(��?��?�����􆑬0	@���cfYZyJ".���?y��������\���lk^���J�*�.]H }B�)�S����~�f��:m�04�#*�M������D�O�6Y�%?��1i��I�Q��X��-($�Z��n�\b��ҝ>���[�B6M��qʊLZ��.������ ���P�6��i�/��Ko��h5�� Q��d�D�_ v��O���ܮR�E��I8�ɓGmʙh�	�o��2<L�3��i�"͓ a6�E4�Ʃv���'��T�Od��y^�M��O �:CB��f	�.���33�wӂ�B;L*�x�(`�Ԃva�?7��m �G���1w.Q{�+h�#g��L��rV敺H"�'UZ B���ժ
]w���'���Od�d��u�V��Û[?|�9�/A�
�R7�'���WoK0��>OR��֟�^wfH7m;��%�)�;K�e��R+I�Lj�'��X���?�/���$�OKr�'����O2�ʗ@�uw��w�ÎZ��}8&%
}�JLQ��'j�H�QB��<A�jnz݅����!~w^1Kዚ�z�.���`֣\�  �f7O��w�'_2���uG��?!��؟���W?�Y�Sk� A�=��I�)>�T�F�5;>��{ԡ̟l���uG�O��B$H���)pӮ�I�
�T�N)"@Es�=�v�ñR��M8Nf��Y���O��$�e�f(�Fb����D�O4M ����O�b)��M�M��,�Ǧ}����#bZ�T"�	����	�?1��<�	�|��EN�*y�H�t�*=���IB��M� Ŏ�(�21X.O��$�O�i�qO���@K�Z�5�g �!b�l��S"Oڕ��[d~�L0S�	��$��ip��'e�ɶ��	�O����|n�!�.d+�荎}2p��6��2J����?�)O.���'�~�L�! L.y:$E�"jJ1��F���'ў�1�1�S��P􂠅E�TK�"O"%�4�پG��S�
��_�� "O��Zu�%j�vxXF(�M�B���"O|��&��ؘ[79��)��"O}Q�N�	f�����+��$�"Om���J��`��ȯ@���s�"O�\�"��t9�|p�k��
|�!"O ���#N�d�B��I�����"O++$:��N]y.�he\�H5!�d�<Nm��#�*&J�����)D��t�Iޟ<��Ο\���6�� Xw�
�>���2Î�j�P2޴�?���?���?���?���?����2H�.�7е�v�U.%��(��i���'�2�'�"�'%��'O�'���"��3�R�p3c� d�R��yӐ���O����OD�d�O���O"���OL����Ud�1+���="@���d_����p��ɟX��̟ ��͟|�	柘`��ӛ�4ꝳ\T�I%C !�Mc��?y��?Q���?)���?y���?��Z7it�Y` �-�\�
�O����'��'�B�'��'""�'�2�C��re�ed۳0�		�G��-��7-�O����O����O����Ot�$�OV�d^.gi�`yu�̏:�r�ƩJ}��m�՟���ϟ@��ß�������(�	+,V�Xr�c)TE����N5<�ڴ�?	���?����?��?Q��?!��C���c��O���! �f�7{\؀ճi���'��'���'��'Q��'�,��LGn�D�Ȕ�źl���ن�zӀ���O|�d�O����Ob�d�OP���O���w��p��Q�@ 	�ƭ�C-˦��Iϟ ����H��ן�Iߟt��՟d�6o�3�\�Q.Տr��=I7���Mۘ'M���Gn[	g��Y�4JUV�)��QMb�(7k�f�<aG��1P�i��T���'�����7��$��ϻu�`kc$�R��Q |�(�����XH2�^�?y�j�5��hWBLBZwZ����dX5��X���k~����ҭ1g,�䑁u����["�R_���rڂ��TbO��y�mK�ɪ�E�+����4DƵ�?�,Or�OJ�@H1j 1O.� ������0=(-���	>>($�G�'r�H�OR�']"�'��!���O��8el�sf@E!v(mV�5��Ǔk�*�'j7-^�fJ�p�)�{��S�xhD��I �F(0��0@���@HJ@!��'���D�O`���������#?@�K)1TԵۀf�;?+ޑ�m@��\j��%X:�r�f�'������d�ڨ{�����F�zI��ׇ 1��B��$8ҭ�>s�ͱ���r��` y�D��4v�<�]5Q��S��O�D�\��Q�ÉZ��A�r펽e��<i���&;F$��+O>�z@��a�ӭV��,��(�f�.Њ�uy�	P�y��O$���Oe��nL]�:<˰�TV>�����R}��'��(
Bǒ�
:O"�kɟ,��3�E�nY�AZ?�P���� m:4�&�$��d-%�x� ��n�2�B�R���Ox%BR�p=��SKP��uka�!� ]��O���Or�d�ORʓ}����b��?q!O�E]n�a��D.y��1�4	P��?���iO������DPW}��k�8Hn�qJl	���=�V���ޕW&0ꆥ]�y������?C�66ÄD����l�7͕�]`��'(�.O�,�� �\/��9�&Z�(a �A#4D���On���P|��c"�i�O�Ѡ�αo��r �/@&� ��O����O�M��	͛oV��O��n��h�/��0��L�)�q�_N�h��76�D��3UB�Dd����W[k���(W!�P�q(�-K�eM�2N�c'ԀEn�	�D�9Y�����Q��p�'0*I
�ěQ�b�'V"��-9�}!&F+t^���N��'w�ɬ71&�����Ɵ��Iޟ,�S�
F�Jթ���M��4��Hgh�˓Y�ǟ�mک;�|��a�f��pݟ`�Sa^�V��$���:1����oϙcje�d����*�'��^�X���ߔ�~�@fl��جH���AB��P�VYQ��'r�CbF5�"�'�R�'��Z�@�ЄA�rT�1��.*@j��ዶO�.@
���L�	��M���>�=�'���o?��n�"����WoIt�,9�	�>c�6��:�$I�$���*� �R9O�9�����uߴ�@L��O������X��ER��\g�Ѽi����}��$(��O����OP�	�D���'1FRy&�̛ 5�`��uG^Ei��
�H�\��Iџ�	�?��4H'���ib�>b���Y�~2�Ō.�7�ݦ�s֦�� �t�Ѥ-�S�mz!�;~���!��z�D�P��!钃ă|qr�:v2u�ɑt갣.O&��ɬ+�x�a`f�՟�B�,�'f��r![ i��l;�؟���͟��Ipy�hܓJEČQ�'���'��9�1&�f�����]%������'�\���Od��'�r��E��e?A��X
s���l+V|y�RN 1'�qp����f��8v
�Xr� ��n-lʧ<��5�	�M���;F�0��+� 9�E$,�����X�	ɟ\H���l��(&?5����\ΓG��y��G3�m�ÆɁ~�Le��P��X�dK��	��M�����'�4ŏ�8�nE����c�:�z�Ο�p؞<R�dV�~��6�Ї$���y�lq��j[�qϓA�Ѣׯd��Y�cZ�����a�Ҵ��/ܵ~c�AWU��@�/.�����W��?y���?��'~Y�X2c���*���K�$�� �f��%���76l!1�'�O����O���͞_���O�p�� &V�<}+UJtYVK��F�˓�?��4[�����Jd���,j@NV8���܊���#�
YJ��aܴbiҬ�'<i��jI�< �������q��A4�B���[4�rj�o��}��Ձ���X�����ޟ��'�D�!�'��~�$���v㶧�5�B�)N�0d�/e���D�(M��ɰ��D��u�۴3X��#%vL^p!�Y#S�2�05,/NJD�%���2�N�̓Q��Bգp�7��:0˧!�����N$�v/���hĨT!#�	��/�R�'���O���a����'�x��v  ���3��Ãl6�Eb��'b�'tdq��Z�R�'��7-�OP�;s�O6!x��-�Qcfb�C�(���'��~�C[���:q�iz��C�*I�N���֝���e�\�Y+�Ԩ�4�K�`����� V�7�aF3��O��$� L@�x���O����O��v��?,�\��˶JT�Ж��O�$�<����=Y�΅k(O��$��=�#A����k��@҈��a/0G��=V���M�w�i���(�''B4�e�	z" j�+0 �cF�Ŕ0��ɳ�!�%)�5;t!�*f;Ph�i�<j2y ���AB>����s���n�����ӲnE����O�?��� �P< ���?���?�����$X��ucV���h�ҩ)�@٢ԍ!�
W�p�d�O�en�����g" ?9�X����4|��a�c�ף\nf�����F,�չitȹS�&ɇ1Ăh�UȆ��y"�֙��䮻 �����!�?����PJR-i�B�/q}�	�"`� ��	�#�MJ������	�� ��+rD��O�  �I�/A��sg?s_�eJ���w������?Y��� ��|���mM��9�f�чb4���5�T,���C�v�P�l�,g����A��h�B���	\"")Dם�<�0�A�j��Igo�U�P��(�?�@CY/g��DKn�є'B��D�
-Ӻ�9���O~�&��H�B���;'��'�O<���O��<i� a7�	K��?i����u`\�!"RT�#�O
͐������')��A��6ld���B��O��H�̓	tl���d��sfȻv���a!L�<)���$�T�u��0N@��O��<j��!����c�N?.����X�B�:�� �=(��$�O����"j�Qj=���OB��y�tb��G�"��!K���L�"ّ� �O��pfA�.n��O =nZß؁%-9?���6�[v�R�y�|PJt�̨<[V}"�a�!n<��$�i�
5�$�G������#t����º�
x��3[�̜�ώ]<�� mS	G���c-O�P��'��BU��L��ɟ���l˰�
�x��Q a�
6;Q���Syr��u:!{�'M�'�4�Q.����'�hE��/K�{U�5a��K~�� δ>���i
�6��5v��סQ{�rʟ�\��>aj�0[4�]�B��$��!,h6-�i��		/L�	w4OH���<�s�'��y3g�4?Ly� C,#����&A�}\�@�'%��'E�'��"4���T,��<� r�K�Ĕ�M�*���jH&!i��'yh7m�O^%Ж�1�O�)o
�MS�+."����K�9��<�/Bj��t���ݢ1;�YR�E�<�&�����ݎbو �RQ>���wV�C�J ��D�E�I����N�ܐ5�O���OT���?z�����$���دTbFh0�G�4��d�O��DB�m�8@����O"�d_�A�	2]V��2_bJ���%�'w?A�a ��$[��O2('�P:h�,6��\a��h��r���<10��C Yۤ*MO��@b�ڥR��mRA�O�ԩ�cTyB��O��k��9e���O����> }�A׻�I��B�H9���?�(OlI[�������?����1�E=D]�D�S��\�L
��C3�`�p/O!�'�7�צ�9�魟��k�3��	S?s�|�XqV-bvB� �%�3(��17E�� h`��WL�-]�	�R��20	��'�8
1g�<1פ�6�=*3$'(��Tզ�6F{Ҥ��'Uj-P�'\��'|2�'���j�ۄ��*ΠR��_�E"Dᣨ��J1�A�I�d�ܴ�?���x~Bb�>��ip`�SBW�V����A�'m��� qDa�L�!�ج��4 d���dDp�b��_�Mҍ@����倾t����ՂA�u�������M+��'��<X�nXF��'���OՐ�ĕ?9{�Ď'�z��@9)2l���L8�lL�e(�O���O��)Q/!��)�OH$lռ��Øw1�|����#Jz��5�W��M3Ѿiݲ��'
.�Ja^p�tc<"��.�0ʾ�Q�L�"&�����1@�
1@�ɟ����(���3Nm@ʓe@�ń�4�4I`P�'$�Q`s��7@�B�'!��$�%�'%B�'P"\�Xط�ԓcr�P���<�ɉL֜�K4��t�N�H��1�&H̓;P�Zq�Ƀ�M��i;���'�P����\_���f�IL��U"ARXN�̓W4ś��`%Z��L��@Z�?I�@�.r�Q�D��@������Q�����@�OF��O�	y� Hd8�����$�O��	q^���ST��y���C�O�����m;��H���O>��˦q�ɓ�����*]�v�2�j�ͧ_����DXip��� @��&i��W���ꓺ�~�aBg��:�o��'��.��Sg~���D,[n
���a	`�J89�����$LƟ�Q2��0�q�Iҟ���?��ᛙgz��F��h -���O�'Ь�'IK	:(���Z��?������C�$�J������U \�&���$;����Ir�8�hS�Od��G�Z2C��T�O��0M�)�b�Y¥�/8�XL�a�� ��X6���y��W�`pU�	�N��)�-O|��� rh�Jp.��Z܊�?V����6V�L���៘�����	DyRm���S<Oe�r$>V�`qV��=8��t��'v�7��O��1r��,I�O�mZ��M�ȁ�%|�`��[�Ok�5���,Æ�X�hM�`��<�훱;��ݯX�BՒ�Q>�`�w�TQP@�y�؃�j-"�>��6O���r����?1��J�?���?Y �SS�f-y��S�SN���0j�!�?9��?���R���p.�d�l埨�'���t��FȄ��P�WoI'��@���:���J�5��(i�b`���-,�8��3��$��a�����˳b��`*g��Epj�P�٬*?���)W��ݖ'L��D�0.�^�C���Op���O�-�%����`�Շ�m�,�M�Oj��<�A*M�T�����?�����Y�/֤�bݿ1T�D@��P��A+O��' 7�˦y!Cd��d��W�T��A[���)ui��R��`ˀ`ё�x`bQ�ߟN�2� ��Հfa�g�)�G�OJ%!g�FgyR�a3�����"��M�p(	x?$�D[�5�Q��M�O��D�O����O�˓�hx�JH�-��q�BA8`D�t��k$����?�'�i�RBT>���Dy�'�L5� L��6�R��V�Q�UО��i� %-D!Y���#���yRa�RN���;,�"�Qԭ�?)�A��xݬ��O��,�֔	�Gg��y�I��
��E�_ܟ �	��S*1�d�O@��a�+,I�ó���.�\P�fG�lA2q�*O����*,R�<���æe�;���q �;&�0�dg���hٴa?���ɼ�~r�c�0�����
aƔ�u�%A��a"��ثK����`�V�>�����O�-hp�
��?���@2M��	"�?P#R���9��x�h��V�3-��URA��co�(����?I��?�/O�i�p��6l�pʓ�?9f��O�t �cD&��7�	z�HM���$�Y}� m� �lM;��	�"0j��DF��[P4z6�լf�j��'`��<#���F ,Z�A8O���"����J,3_x��%�" 0�i	A�R.�K�C����O�D�KPU�N=���O�x��;uc�2>����˕�g=0�V�O@���N�w=T�d�O �o� �fc=?��'T�&���D� >A����*��D�hՊV��n�B�r �i�^�J�fDm��n�@��p�	�l)P����q0���$xԭچNG�t�]�J�'�Dl3,O,���*Y�|�z��ן�I��������Y��@�	#�q�5�X�hj��b��Ty�R�X0e
��'P��'��$���$�'��� $(<e�E ��(��ģ<����M+e)Kg?	QO,��L��?a�&%��%� ��`JA��x۬H��jj����E1O���S�%�?ن ��#剶�?Y�W*� q��{<i��P��|YS�kS��?���?i��?�-O��bU�2�,�D�rHA8$ #`8�f�́���������I:��T�I�M+V�i��R���;	6i�'M�W㌙9�T��X{b+ֵS�k�l���B���,��.�L i�(��]�;L�к�ڸ'D��4(��g涠2e`U-p:� �	��`�	�?Yʃs�����s!��4X�9҈Pm$8 ���[�X�Iߟt����,�l��ş ��4�?�A,�t?��KO1��}��e�;�ڵ��L:Y*&e�P� �"�]�M�'Ȉ�BZw�x��Ⅰ}fڙc�Ģ]�Nh�"�:)2��_
�5ZU*ą%Zlk���8��>`��rd���,�	��X �,JnI4X�S׉�ǟ���Xy�Xr�$��'d"�'P�DI˙tsʍ�R���dxa���SN��'�<R��,t�!ߴ#�F��DXx�H6#�?B$fEY^������W�x�ᑬ!	b�x�'Ȏ'�ؚr;O��]�+�����'	M�/O�X�Eȭ�P�@Q+�B<y�l������
YWd��Iߟ(�I����	By��,� ���%U�#E%��C	
$�V
?Or�'`�7��O\��"��tI/OP�D�1K]��р��\UЬ `�:�7�?R�X9UME�(2��{>O���)�uߴ;�6�O��0+�X�Mx��m���Yٴ�V���9��'��'?�Ĩ��v��S;H|x�G���x�V�����wB% "h��O��$�*�[T�?5��4�y��4
{���#n�Y@ףX1V=�f�c�X���OL�@B��)9k��݂J��1QOO	?����Z�{����R��?)a�W/ey��I�o�y�'B��d�0i����uD�O:������|{㭙&�E����O��d�O��$�<1w��/�6q���?Q�jAz�Y����#ے�)��:�u������'��=��v{ӎe"�O��w`�zM�́%H�3^J��×i�%���[�'���Hظ]	���'�Ց��i+c�"�PN�4��K/��)�b�ڒ;Ƥ����4�����0�G�A��'?�I��Tϓ
R�PR��a/���.Z'����	�2rHQ̎�p�I��M+�PH�'p�T@	 -�Lh:t(�,�Z��M�%(ɦH��@Bsm�,�ؗ�#M��%i�d̓I�Rd#6Dr�7m�!eN�1&��@{l�Q�"֧=�H�b�<I��'�"1�0-F�`r�'d��Oϔ����2�X�%��{�J�uI5k��I<x�aZb)S� ��ϟ��+��S�<8A��0�����*	4�����)���������4=n���Q�(��'`�5�t�"��;�����Pt|9)���H�bn��u'�Ot!b���Iy"�w�\r �M+ <��a�/*�LX3C�5?0�){$N�O���O�D�O<�7<P�J�-�?� b1�*�j$�Τ��E�b���?��i�R
���Mw}RLt�>�l�"������+w�H�A�"u[(ȑ�ZiF"iӂ�)9���	��]�$����4�����ݼ��gQ[�d�B��(���q� ��9��B쟀�Iޟ���Xp�d&?�	PZ~�x�bB�DRj�W�Z%G2L�'|"��%	���p�'$�dsӬ�ċ�#��D�l��2����\�"cK\ 5�9�'�n��Sr� �4���N��u�o_�vO�Ă)}�~$�w�>rGdH��KڍIz��pCB�?Yg.O�O��	2�?�W@�<|�����?���
��Y*$�C  ��I��
=M@������?�+OR��Ůʇ�F˓�?��'�Pi9fȤuT�T����)L^p4y4��$��$Zy�'c���
�~򢂾(�ܐ�'{ĔxPOY�"�z��#t��<Q�d��cB��POG$�IҺ�Ufҟ���-T���DIc�,��DH\";~5�D`�?���ɻ��Yb¨���p��ϟ\�I�H�'�鲐�ӶFޘ���$�2\žU���F�c�RC��'LB�yӶ�ĉ�&�I�����ɦq��a\> �|� ��S��#�l���M[���rE[���27�l�Γ'�(�$�j�e	�#Ψ	a�)��u��`H�ƞ1fe�����rz�F!��,�U�#�O���44z����5L�$I�O�<��
�*c�l�A
�(!"�L�e�����VK-�h�r��ɯD��]�A� w�<��	�&=�������HY*���	a%J�r�.�
�Y @�hm2��#)-Ƞ�"q/Ց4Lpj��u�>r��`��7���� Fl�x�1j�8��'N^&g�n�r2Aذ�?�b���jm"0e@����?PB�H�M�	��R�d������𰥍
���P��ן����D�'^�	G}2GڊK$��`ʰ4pе[G�T&`s���ѐv�Q��E.>m��ںXH���+��lP�M�)�e��(ٶW��C�ɬj�:�$�*-��M��ʄ]�J��$�%�^}i�n�=
^>�ʥj�i� Y2�b��2"j�/k*����E�;������+5�ά��'�%Vp���N�Vm�o�55�,�!�J������L�3NZ���F�9�X pn�����X�pQ��P� 
��D��Lߖ�d!�t��7^H�Q�� 9����V��,�T�=1:%�R�Z��򤘷t"��'9ɟF�$�O�\��*ϭ.�ZI�C*C*�H�(E���d�<����?���$D�/�����5��RǨPq)�%�Rd��;�,�I�k��d�O4l;g��|"��?�ި�?i�K/F��feJ�Ed$������$�Od�D�O˓B���s���h|S����C�Y����dG��d�OJu�O2���'��b1OH�)gHG�b`,!2DI;d� �'�R�'B�0�l�ɩ���O(���d��T��D�\��ĖP��ux`�O08h��'!2�O`��'8�R�Б!�Q� ��Iy}��R�G����	��,�	�0�Lc��-^#��I��V<�'���Je�lm�̗7E�D� ���G<�I�QC 5�I����}yʟ~���J$o�����W�yւ�Y���OhI�@�a��ӟ����?���O��1�0O�Y�'�)�����R슋aD+�?��-���?���?	(O����<�I0[� ѵ)ĻC��;P���CJ��ݴ�?q���?Iڴl˓4���	ʟ pf�ܙ����$J��7$���&g͒��I{�	I4t$?���ß����d��]�R��G�z���m� 'Q4���՟䱄o����d��y��'�r��ɟ��Ej1����.W.����A�<1D����?.O|���O�D�<a��7]�\�x�'�ZЈ\�E�'E �L�\�� ���O��d��|���ퟨ��X�t9����a���S`��#�a��J�ӟ8�'�2�'z�T���sM���㡇6C m: 2;�Qh�/D��P��f���Ɂ(U��I�?i�'��=��4{���7-�֨Y�ٵt�Z�X��'7��'���'�R�'�����r����x�ře�'7U���O��r�2��OL�D�:k'��К���y�'�?9��?a�Z0�����&�;K�4�QJ���?��?���?Qe��D��s�����?���醽l�l�S�h߃$�ne�Ǯ�7X�I�.��c��I�O��d�O�{�*g��<U��x 3%�)������?A��\S ��'�i��O"�$!�<�4b��8����4Z ���*B#gx@4�'CDIsq�'�ʟ�?1� Z}��� 7�\� A*��n�z��'��J��'�B�'l��O�剛Rq瓳�B�Rs��_�LI1��A�z�l�%�X����y(�(��Б�ÂW7�]HG-׬L3b�'s��'��p�#S���w>�ΓH:�
Δ6.6�m� �c�t:��D�	My2�$�O~�"x�|	'$�F-
���ǌ~Fr�D�O��� ��<!���|��'���~i+1���b��R��w0)9���O�ʓ��'��S�8�IU}�h(d.��l�Bi0�,�ZO����Fy��/L|"0OT������y�O@.D5�W�� �S� ,�?ى��'	�������N@�|���Z�l2�%�$}��e	�f��|I��	�Hϓ(n���*��|R�'���K��0�Zx@��<���?y����D��XL%>�� �@,:#`�S$m��2���(G������>�r���
d~��|r��?�'*�D! M��Fs0S#l�AtL��ݟ8�'Ri�5WP����X�����RjB�/����J�i��}3`�_�|������${���-�Ļ<i�dݽiڵ3VL�;mj��C"�?�)O�E.�ܦ�O���O��ʓ
Ζ�BրC͞}q��X/1��� �O�ꟴ�I`*I�	����Ky�[>��
���M2�%Gnx !� E�w�NA0���!JP�8x���˺#��Y�Q�����b�І&3��bB�5H��݉i�XԲ��'�'�'%�N��H"�'D!;�BB�V��@B���+��' �'���y�=�MÀO9I��F�Z8Mt����'����>�O��9O����O�)@a�x�Ȭ��,D�O�%�(,��6���X��J�	$i��mk"f�������xΨ|���x9��Iڟ<�IU�i>�s�Ƣ?��s�P)Al�]Y���+����S��On��;��OmHu�9O
�����R�1�@Å3,�4��m�O��e���Eן��o��	DyB�O�����d�?�� �F�;{W6dڱ>O�b"�'���O�.h�U�Ů��ܩ��'F��qV���W4��4Å�@�F�m�򩘅"N4C'tx���<v`��0ת��C��S����0��ǧy�~�!rK�"{��1%$C�P�lRhZ(��XR���YVi�I�-��ea�I�(o��\�'D�L����ߓ=�T,z�L9{��)ǏB� 	�ɨQ���-�O����O���Ɠn� a,�OL�$�:k�(!a��b�)s蚶E=J�ʔ	\/�q9T�>�O��x�/E�>�tzF厧`�� H�; ٌ|���Q=�+Gdm<����*r��'A��Mw�%[��D*1��@�'Lf7m���5�	MyB�'۱O�Aj�`�i��E��ݦe],�����h�y�O�X�I�B>�N5�$E�W���A�%�$�
m�b��<�2) +�ђ��Ms�`G(��8��H8F����ӎ���OF�r��°iJ��d>���	�q���S�J�>9��+d��0�U˞�z�T�H�jUFX���Q-�$�D)@c�>�a)ҝ:i@�F�M�1B��3dDX��b�I�O80lZ�M��4DX�!b�hΠ/L�C�^/Q�@�U� �	S�S�'d1>��ٖ~��q����^��?ɦ�~rNZ%{�.��&a�M�\�b#�C3c!xH����(宁���O���|���M�We�lf��� G�p����!��_��'�hk���d M�O��I;�d֜S�*5�ԂH'B��a�'	Z����i݊��Y�E(�>� ��A�G�'z��0������O?�0�SO�
e�<-HSj׽gNx���'f� "� ҇.N����L�:�L)��	\z��h�� �^	:Q"W_�rLp��&s��r��6o$��'�ȟ ̐����'���'oK�7�~��'���6=�e��Q��:F�׫��	6{��	Di��n�ў����Öe����G(��~�T���; ����O	����e�g�	lT�����*'.=hr"7�.� ���?���%&\s�S�gyb�i��m��L�X�B3섹1.�y�?$�	9C�ʂ��sN�����O���S'��Gx������Ic}"�؁$�B�1� �8?:�q��?6b"�ͼ^�0�$�O^�$�OhT�EX���O M�W�W�3"ؘyա�������+<U3�$���>94Ɣv��D晩.R�!AÔ?��!�j�%k�`�)f4�``�I�V�h�1d��:٬�q��ˑ2y���Om�$�M�����O@c�H��5*�M��L�/�d#u�%�I֟��=A��|���<锅qb�Vmb�(��M=d�DO٦��ɝI,��ߴ�䧯M����k0��k|�z'ش���'nEj�<A���f��t��0a�B�XԮi�� ��Y(3�S��пy�����F�W ֨C��2O��!�"O����G�4Ϧ,�w'͘R�ֽ�3"O�Hzƣʛ[oF��O'D��}�"O��@u/G@��	X�,��L�"O�T�񍛂0"0�)�l���"O��+�g�1]d��9�C�W��a�"O� hU	q*��$�6ı$��h��X��"OL�{�L��5�J�{����"O.�C�Ǽz�`}�B�J� �6l8�"O��[PF{��R�����("OcA�ķY��9& U�l�p�I�"OH\K (���|JҪ�GQdĻ&"O\|�4�Z)[�MC�'��*E"OJ�ڗ"ƯWjν3@��@��С"O��������I�E��v���P�"ORԣdɍ�.�،������"O|���$�@��Ua�u� %"O�����/���:��և$b�P�"OVx��oϲ"��Ƙ�zA�0	�"OX���P�
-\�d��`ã"OV��í�5�t��lĈ@X#`"OR	��D�]�F����.����"O4B&�^�N`�Ӈ�Y	|6"O)�ǨC�w]lI/e2�J�䂫�y���tdC֌��X��,���y��q�jC�3z����W���y��6s�|�ӣa0pV�ݷ�yn
&:Q���UC�xA~i�B�X��y.GgNɻ�KY�	�6A�`� �yr��
�t���@"2ep�����y��ܻiLF��5�ƈz�����y�A� ($���6(���O��yRA�$#��K�I*"R�`�� ��y��h� [f�\���d���y�o B7�qW{56�a���y��	b-�����,i+���yI�	z�!��A�lvȨ��+͡�yb.Ș`2��Ơ�?K��}:O��y�D�)4>��c�Զv{�B�(�yri}-�dȃG�[�6�8Pc
��y��Ǔ!�
� �L�C#�)��Y��yRIU�2ֺM�A�:vfY�m�yr.�)K����V��N#$Ia#'�y�IֱS�PW���@H�d���yr�O NS,@{�������@*��y��\�(�,��F���|\dG��6�y�`���(���E�X n�9�'�%�y��dL������+��D�����y�o�i��q(C� K�m�G��yB��%jxR��J�>S��02 ���ybI\�
����k"S�p`֞�y2��	k�x�zR΂�&�2���ր�Py�'��=����k����A�h�B�<9m��u��T��M��+�Ay1�U�<!v(��.�`V	<l<>���z�<���O�H�^y��d��-z�I�~�<�cfĶ{���S)[�S*h���6=gDh��?�)��<�'��3h��i��ͻm(f����l�<!����22��A.��<��t�!�ꦕBw&"0�m���'�Tx@�k��7��H��H�Sq\�ӓtr�E�F$Ψ:*����25�p�(g߬0s�0�GK��	.tZ�)��_�1� ����dϰn�4���K�� ��J;��'��,���O����V,aN�υA`ބa��	�3B�� Z.v,��4�ȶ[�&4;ԮY0N	��'�p<Y����g�	1��w��%�J�v�ur&��G��![&� Q��^&c����s��UJ��� �$7A���$f�-��Y1J�QH<��"c��8��t�,�Kd�04f-�f�J�X�˒�Ga��@C"`��5xFw�&�SD�Y�10vM]�X ���b.��B/}�~�c��'S�U�'R��`� G$;�F Ag	)V�����A�=W$�av�]�vҚ�R�ꋩ>�s��e��)QWmɩW����}���`|B� ���(�a#B� ���n"I*Cf�-�)ەlϩ�X4�6$3oB�: �2]ɜ�a��Z ��HAd�J����ʘ�U�%��
�F�v���S�?  ��F���)�A���{9\ J�:k�"��2����p����$���6�Ҫ,�e��4 XP�4q��*7/�t�:9	G��)�Z{��<����)��t�n$R6 GD���S@ҹ�Vy:�.� `z�Aԉ�-78����T$�M3T��0�,��u&��p;����ݳhPR��#G��:u�Q�@h���d��T@�d	Ǟk���r�ZV�Hłv*��5 �9�4\�u��]���U�i�XQ3�Y��M�q��.��\�^���@2C�1O�I��*�9q~�U�F�'{�P`���>��NL�ȍ�揀6/�HE
w��������܋o� p��T�S1��q��UP4����[�l��Z��ق
d����:Y�����_�a�:��#�4 t�@�2�MP��z�(�;�PQ30G	&/��@� 垯e�,А�ȕ�x�xҲ,L^��f�w��%�d��\B:[u
M,���^;M����m�':��M	�Nއ8���
S��>�Bu��ٕ#��I�)O�0�=�3��%?��iIҮ^�<���j�o��v����RA���
���&�(9�	˓3�~)Y��%]G>u2�;=���pŔ�5��@#�@�=<<�Ѓ�
GVD	{����18��@6����23��8 ��O��v��U)�C�"������$�E��!�A���) zDA�27�D�ȁ�ܱ�̩�R朠R,x�P�H�)��a*̏Mn�)zu�
0�����.Ѿ�����b}�/4-�����]?��$Т	ShE�R�ܒ*gН�cˀI�ڀ��)��-�2f\�:�
 ��Q�\p}���Z?����)N��
4���}�������	 ٰ<��c�:�Խ�D#P��836DM�������H70p0E�1fN��*qj��<�ʍ��cU��$FD�����SL�w��M1%j�-]�i �5s�����T��|TYa�(���Zf]9w۪��Z�dw≈*]$g��r�mJ}@��9�G^
m�ȍ8���.1Ӹ���d�`�ئ�|���쪡9�d�2O�:eѴ�T�>��D�Oy�򉟫vp)�� �71�xb���)�⽊�g֓-	�a3��H0,td�&#٩����B	�f�(��%k9����O/�B���J�V�P�
�%�R/�I���8��E�T.P2�	���_�Q#ʩR�D�ja�W$�}��A4��r�m��X�E[�D��&eε�r!9b���ā�[���Lׂjk�XH� ��^sP�9,]��`��Ɖtؘ�էDu��1oZ-���0����0e1�
 "ݾZD�);��<c�n���'�l���E�N�����oM����T���{�Ra�$j�]�#�L*���Iuӎقb̼~V\I"	D�_�4�����Q�c�,����+�����كa�D�O��1k���	���'=���jP�л�-c ��K�ty�[�q����mU$�pHy�@\�=X�I[�hʬU�ZQb!O�T���+���F��q�#ԕ䠉cĩ�9���"�ښ8DUYPZ9E����+��A��A��᪁c��;�5�D�/9�n��kN(�KD<5F�B�/8�y��R���*�E�F{l<�"���>�Q1��/\��R�GƂ+���Q��S�����ͬGzn8�2ϛ���b0� �f�~�d�Z�� ��<�V� |�h�bd T�p
��jP�J%s�H�%�<Z�� @D��:h��@��T>Q�<��%IFpР�F�
�s�J�5��G�w� ӗ��f����N	6j��'����I�h�v�Rg��2|�O���p�.t,a�ƅɁ{�*�K!��!k�]X���&m_����'n��B%�

<C�aG⓯3�,ls�F�-V����D�v%<�:��B���4�J�<B���'f<˓,�\�@.�7+2T��֣��uژ��ȓ��4uo�1+���тAʊT� �o�'��!*V���?Q�j;?I��(x��O�41f$E) ^��w �oL2��v�'h�xk���w?��,��x�x��"�!Ҕ��v�l�	�<Y��8�IB�J7@����k�¼+�㝄(��	$%�Q�Xy4�&"�d�j ̈́�X�4�CJ#D�����!/�� a��`^��kF5D�T呗u���)]5%b�cB�0D�(y�@la
���Q�p �Pn(�(@9�D �:��43��%hL�"UmۜB6n5��Xx��+p�E� 
�a��Ù'�Z���'<K�V�F�mP�p�T� q%�#Lx%��H�'��=9Ҥ7�U�?[�ۆ	�-/�M��$��Si!�$�O������/8���#Q�E�!��ͣi��)�C�	/�3��/{�!�T&��ہnW
a���v`����'��Dy����垔!��H�x���#[0�y2�,("N%k��Zp.L�D�V�O��"Ǔ h���+��f8���țO®�ȓIWj���D���|�FE~�����Qa�ݾ8� ��$[�H�D�`�jT��y���,k��1 4�ŇK�Fe��e��y��Ce��"�C�F5^]�[��yBE} ����H���R��8�yB�I \���Ã7E�P�!�J���yR�B���%���>���x�����yr���W?�t�F璆?�B5����y�N�:o�Jt���X9+wx��Ci��y
� @��P`�
ft���S$���"OJ��L�.�@X׫R�YIFT9�"O���Cv\�YT웸K.��"OV|cG�P5]�8�놜Y=TDC�"O���CD]D�9P�E#�E�u"O�\��$��p�U*��j*P9��"Ov��R�Y<1Y�]"	V�>�aJ@"O\-)D��MlP���L������"OL双&��Q0«Ѥ��HX�"O��%��"!�T���J[�����@"OL�36+S:W"�l
(֋fa�Z�"O�aj㋨V�ąs`9k���"O��Q`��	F�K�Jz��"OxCi����U34�[6 ��!"O�ժ��A�V�x�N0�b"O�����u� �C!�>O�p��"O����6329��b��?�nt��"O�EQ-A35*�g� 3�4Xq"O<� �F!J�^�b�,�4#U"O)��ԥ.��DS�����yi�\��#�o�3�ઓH�y�۬I�h!��푎/B�Xy@
��y�h�pl~!c"
���C��y�n(;��8c�*Q���!K��y�=,@L�sR�'-��E(�y��;~�Ȭ�3i_�� R`CO��y�	*E�ZU��`�.�Њ ���y��ʡY���� m��2˖�á�M�y��gʸ	; �܊Cn��q!H>�yb-͟)8l�U�̌Lݲ�{�@ݏ�y2��_����`J�S��µ	��y��
����P�p�0�)�Y��y"+�,j�p�B�%w���QV(��y¬��i6����0e��9Q5�̀�yR�J+/�l�V%��gI������yr�L'� e*XN�H+H�9�y�I�=��y8G��
\0'����y��[�&��B���(xQ�aJ����ybHL�`8m#��<eR��6�(�yBۥx۸��čO���@ƈ���y2�D���f��AH��B� �y�յWUfPQd׉EVb�x�͚�y�N\�u�R�%��؋Њ���yr�D5��B����7vp���-�y����M�4��e��,����@B*�y)<W��(��G p�h�b!�yr�yf��!!�Mr�,��Eb��y���07�������?i���t�H�y�r���)
��m�c���Py�&B"cSR@���4�A�f_z�<��d4&�P�˔N	��ޜ#ᆒ^�<��FĂvm܁��jS �4�k�/�Y�<�+�b�M�"ľ7��<���[�<y�C�`,4[ь�;v��$
�M�T�<��m^�U��$B�R�r� ���)�K�<�a�E�4�v�B���K�49��J�<���� qf̋$���>�JŰeoM�<Q��Dt*��qdS�efl��C@�p�<�Ç#z��lWdU�,�4Q���e�<�k�*A�+'���4h^]��,ZI�<A�L_�f�|"&O�`6�p bÌA�<Efǖ]���%[F�(ɛ�L�x��\�&`��M�x �Ю�TⰓ%�ރ&Q�x���ӡa�,@z�"Oz<c��
:��"����!�4��E"O� �u��N�gz��@5C�.�&�0S"OJ�p�$��N���b+�d�J5�W"OR��5���6�����O,qҊ�P�"OH��4`.QE���#□$�Z�1`"O�tj2*�3h�l"�A�1�D�B"Opa*%�];u�fq�5�K�g"
�)4"O�t�����+[!CB��K�Z}R#"O��&��'��i�ң�al i W"OJ4�����G
���aM�XtH�q"O0�G�˂,����<���"O��J���K^�(Q28R����"Ote��� c@��vBM������"O����L�g�n���]<��@Q�"Ox�{U�ˇ) ��r�	-v�����"O�!:�-�{e�N��Uʧ"O�%g��#!tz-��A ��5Ig"OR$��C�I�i�2B��G�)�D"O�${wE��o�$Y��o2{�b��G"O�hR�̍4"�\Po�	'	ZX�"O:ࡦe˱{+���+�Da�"Ot�J�bؠ/E�����A�|�6 @"O��A�[5,?Xi�Kة6���Q"O���g[������C4���,�yr%��1��x3��W�E���c2G���y2��h�*�I�I��l(Ve���P��y2���w�����$TLn���%���y����T�9$�7Gu��2�#֝�y���@IV��j���`��y��Π(��0G�¥/��Ha�c��yBg������fI�&�((P���y�Q�*�Q����
S�:)36hG��y�e�1)��g��Q�U��jX0�yjXD�:vF]>��E"5c���y"���}��P�#j��0��i��B��y�CQ>r|�ؓ��+
	��� ��y"�&���xӂNS�<�#�
��yb$Y�^�@}Kv��!D���R��˒�y��Ygfd��i��4q��k#!B�y�IG�.�ђ���'�\� �� �yҢ�3._(x��ſPk����y\>Z�
mH���=�t�2�J�yb�̲f(y��ü6nr������y!���=�� U.�ҁ	¦���y�D> ��E�6`ŝqZȝK����y���rOj�ԡ� ��Yp�ԓ�y�o�����R�*��q�',���y���KU���E�����S�'��y��J7��a�5�IP�C��)�y�M$Ǯ�2vV.v�RK���yr��.�,��e��m���jS��y�O4K�̄3�O��Ȳ!ֲ�y@�'H�<4�t�Nv��p�1G^/�y"�޿[.Z�S�s4�IȆ����yʛ	!˼U�7 �*�%Af�M��y"C�-�l-CJ
N�re��c�<�L�6�-C��G<G 1I��M�<���
�mU����:9��)g�R�<Q�X���6a��[�&�`nLX�<�$%wX-h���	T0ics��~�<����96�Yd��=LY�U��z�<��l���L6"��f\JA;W��w�<��iI�L��
&o#t���N�<a��E�뺱�'���Ƹ3�%JL�<i��ʄbW��cF��VxL�x���p�S��h��)� l����;!V�P�����Q�vOl� �O�F^8��@lMb�E2�I׬E�X�ēW��rk�68�@�S$!�D~"��������d@
�_A��CUH��
D
(��I��y�o���!�T�	,�|���q	�'�-(�k��ēHa��:-�I�h>0�3��[w>���*�X� C�ɺ]�Ȱ����В�5$�˓�y��OH}Y�S?1#D�i�r ��[?1i�^�6@TE��,뼁�R5�O�P+��Q�_�*�N�W�N�1�Jڨ^A�ո�i��hC�')���S
)#zSS�^$�y2� y�`�JU�,~�u�)Ee�'��qLxhR��=$� 8���k��X���i�;���M#^(��F�Mn�	� ^�HO�i�C�зT���ð�٬���c�'�|I�d�l�̹���P�^h�E�ȇ�����Ɍ[��	gy��Az����T�fI��X�`�u��G;ziH�f�TX�Lb#�?c��`+B��{����C��Vb��0pm�4� �uȇ�4�M`'���DW��r�wI�QMS7O&��"��R?O1��
�>b}�*ѱ�.�q��!HSLp��K
9��m����7���6��ao:��)Oܱxf�$s����N%۰��2�i�$i�D���I���w��`��$�+&$j�H�mn4J���1|�"�c�Dڠ���2�W�y���IL��<R��@�OB�qso^� �$�&���t��IG6��5�ފPuNTRW
^�E4��q`�K0�l�S�\e`XB/R-'�8�3�Ϊ�NUPSN������Y
>���o�?��A�+� {��h���C>FH����Y�V���k	�呠ᘊ/B
26@��O�����D[)Z�� �X0CC�X�O��I��yW��f���x���,G� aCbT%�0>��P#*p*�JR+Ω#��T�?��њAD��s I#��*B-�E�A(���	Z����@:��Rv )d�7��3YUP��Չc<�s�*\�zC���WgX''2*��!����s�T�CT�,٨� u�ŘJ�(A��g}B���~"�1>���([V�'z��.I<|� WM�k�F�aE�/}Tx!^�Z�� ��ұ���L������!��6V��Y�kɀO�*��&�ɪY�~maq�X���>�@%тM�x,cѪ��b���Nԛ�!o?	�}��U�"�E��&S��.�t���e�.)ȉ��ΚY�a|BF�E���`��A�tJ���~6E9�K��'�洫�'L�	��͙צ�R�F{��I�D$li�C��7c���\��(O�D���Y�O�$mk�K��w��O�(����1R�	Z��"��+��N�\L��I�3�l�0�؀[L�TC�)�&$;���&N�����Xd�c�S�,O��OJZ��ߊH؄��h�g~$q��"Of�E���{Y�(A�'�1��IQ�iV@��_~?Q���۸6m��`1,��*P<v���9 @3X��i*`(>�B�9A��U�4���y�D�ş>��[?$
#?!�%�G\xL:��3f�^5��`�O8�p�5ီL�x�O@�(C�V��@�S��Q%ZM�Pq㇭rDl�:��1���Ea�F���@�T6a��$�#��	�^�'�l�S⓺K��q��@gPKwmƼH6bB��(4�p �〦c���+eꂃybj�O��)a⒣����O���1��2�<�d�E��z	�'�Ɓ{`��4@`�����N�mHug,�I�26���O�`Iai�b޼��%Ǭ6����O,�'o�5p-�hX��E�4@�4(�!?rv]�Z���sb՛Gp&L����"!\4���x�&�&�h�F�F��l�%
� rz��;��#D�8��c�5/�иt*K�mvth��+D��,�|�ڌ�d�S�"����a�(D�Ēg�5l)����cS3}��M��"D��Z�H>^�R,�E��&`�6�!D��3�����v0P�Qw�8�ku/?D���%B�-y��rF �L�1%�2D����BI�v nhaqk�
y(@
.D� ����+C��p�(O#{̠��f*D�;�$f�h`�i��fRykq�"D��8��M?�~m����r�*1ru
!D�@b���WZ�% �I\�ux��`!D��B�*�2V�a�@��=g��,��'?T����ꋆu^�c�ȰGq�9�v"OlM# !]�b�����ϛ!eFp�"O�ʠ%R-z�,����-Z|��"On�qc�#�0P��(��'IT%�B"O� ����f��A��<22�Z71�J`�S"Oz��!̋1,h�(��yoZ��"OXTЇaQ SªTXc'R�m���c"O��x��Z�G�Tz��O�h��HAc"Ou��Eݒ~lʈA7oF�	��%k"O���5?Z��`�p(��"O�Y9�B�*$���ʴRk�"O<�JGo'Z0dt��G�<`d59�"O`5��oڇQ,��Y�RQ�}��"O�Yae��,Z�`R���o:�b�"O�%���ߟ1�Va��FہD��%��"O��5�ϙ�`e��G;"��Y��"O2(��.PLĐH�愿u��q"O`y"��Zǆ����47&H�8�"O�I���J.���*�
FEb<f"O8��a���5Z�"�Q7"Oh�X7��d����1LW$�K`"O��w�×!�V���'~VLY�4"O���4]����h�R���#"O&�&w����F�V���hC�ъ�yR�Ӑ $�Ч;�t�q�=�y�"�� �5Xņ�1�t��c�ü�yB���-ܐ���):e�U����y�ń��r�B�$]�"�Ή�g��y�@GAE+�E ���㲡_�ybFA�t�|`�!�@,DhR�%k��y"fG�+��H@�R��h��ず�y��8(���i�S�\�f�;�]��y��0	)�X�O�>i���C�վ�yB��h�n�c���-`֝ҢD�y��Н?RX�Qd߄'p���"�ճ�y�@ĳ-���RR`�������@��y���<��,N� ���0�T��y2G0+٨�`�F�2���;׎��y��
n��XG��#�H\��ܖ�y�A0���삼�&���C=�yR�}�M��FE�t�,U���y�+~��R�ꍴo�8 +�E�y�$$w�"'Ɋ�xX
��&��z�'W.Qp��Ā'����VnW)kM���
�'��9���������C]6��y�_2�$�؆�\*&x����B �y"�� �UPw��/n���K��F��y�č�p00�o_�B��H���y2CE� 52a)�i;�3AN
��yB�V��e�+^�+ M^;�y¯�	qy��p��?T��`������y��M���<
&�LKIt�+�'���yRc� 3�ȑfgȻ9�� F�H��y�@�.b��vn /q�8(���N�!�DH�x)��r��uZԉ0S���Z�!��U�%l]����mA�ز)�">�!�d� ���T�&a$L8ghV�r�!�D�iɪDE�). 	�0G�!��PC��ˠ��):h��)�!�dW�E����ID*���7ę�K�!�� �6��n[6#^1�RB�>P!�֊C��A �L�O��!1��x!��ٟ�~��$F�/[��@�/[!�d�!��B�Ne9`�A� �X!�d� &���&���W7��h� �>wH!��ֶ��oИLz��Ȃ�@�O3!��A�{��uY�M,0d��O� }B!��+w(.�y!��H�Mٵ���hB!�� ��1U�Ȓp=<��Sd85�$U"O8i����0�ŹSW�qV���"Of����%]{��D�Ϝ%bԌ�R"OVUӇT�}���p�G�E�qu"O�4QO@�ffREp#��+ q�$"O։kU��^!��k@�+?�e�"O|�(���,�0��Ҽm�X���"O�e`4�? \��3�C�?>(^�Bb"O���'.ܖ6oD���@5� I�"O��8�>= �yе�G�����"Oy���0TH�I��M��Ъ"OV�
��y����%��~�B6"O��S��g��	��m� ��,��"O�X��`�e�,�:�'}���#"Of���בG��h�&	��Gǖ�Q"O1�B�:���#XY�p��"O���/^g�ZIc�)Z�mG�}��"O�`���G��W�
9`��"O ,X�틛 )vm� lG�jK���g"O�4[��t)��W�X��x�<�Oάp枱��72�h����w�<yg�� "@R����Z�G-H@%D���J�1F����.�},)(��7D���'K�,W^\�e��}��xa�2D�\�����j����`
V;Y+�\��2D�Xc�/HK,<i�A�Do�� ,/D�����?/�d 3m�*�n�Qo?D�|�!-��rf��g��*�l��5$(D�̺���$�is�R��.\B�b"D�t
�f�Q��:�gg�����>D���ξU��AJ�
� rǊ5S�o9D��� n��a*� �W���&=�E8u6D�����@.Y���P$ J�T`t)���4D�j4��V�z�C�e�F�f�U�'D���#��)�
qkɄ�s;�$���%D��#��>Vh��PVj�)r��YdD%D��[�h@�cd]r ��	,�$���&D��C & ��mQ��N �,�`&?D�H:��"U��Ц��
/�*e� +=D�xF�a.DI�����i���ҏ;D���Ł�le.����R3��%:D�T#��P�ޥZ�bL�=��t3�.8D�� ���|�䄺���e���k#D�8#�jNP�US�&�!3Y�"�#D�h��?;�xp�� �H��`,D�2g�ƣv$�y�hռis3d(D�X���3A.��S���,՞��E;D�(P4/��0�� ��]�b�f��b�7D���񏈌u@݃7 ���0�i��5D�$�WJ�6�̡��Ș�t2Q!��0D�T)�C�g0��
X�!��,�t�2D���#Fĕ���!ET���$K�E2D����ޝp�
�#%S	G��G�-D�8(�A����W�дV��@�!*D���ĉ� O�T��J��ez�S�)+D��q��
(w��k�̒}���'D���c���l�� 2d ����ز00D��S�!Z=6�@e�3	���(f.D��8`ϐ?(�fa��5¦�1�J*D�tp@T�$. �!1&�"�@B�O#D�,�#&�VSD��uGK l�^���E>D���'�N2"蹲�G4�F,� +>D��a᧍k�Z43RC�+c�j��v�9D��j�%%#|HACV���c.|����;D�� B}96�M�-�JA8!79�r"O�% �Byt���j��=����"O<\C�
�Lb�f���� 8E"O@�9��-]�b�$(A�O�PD"O4�` �z�� ���+C����""O�c��/Q������?&��<	"O���*J!y�ȽH���M�v�ñ"O��0��E�o� A�a%�bԸ�"Ov��Ř�f���	�CSdn���d"O陁��*9G���7�13��)+�"O�`����$��U�i�)a"OIɦ��g����(=d.��"O�h�dbSf��x��Ŧ\P���"Oi��h�!K�&\�rj��C"Op`#ľU�`�'��x��0"OX1���
"���U�N�-s���"Onݣ���)j�@�v(�(�H��"O���$$R�H���d�>����"O؀z���~�F��G���{�$��"OJx��	�g"���ãJ��"O޽�`�}6B!�t�J z���'W�'��p$NȄ->�`���|70���'8L��銿4/:A�և�
oZR� �'R�֨�D���a��P�4���	�'�����o@�&�V$ &�͌*�
\q�'���a��$c�pxP%!&P�V �'��E[��C% t�(����X���
�'�~!K��A�{0`�;Q'����'k&��w��}F��g�^��,D��'<����k��!���Ɗ���'�^�p�'KH|����:ۘE��'��d񴃍(1��AI �|j�M��'�`���+��yQe��wZ�J�'1��ȗΌ�A�$
��_����'�N�C��Ȃnv������G��'#���QN9ӆq�sd@6H���0�'W�X�ȣ(e:5Aci�Dny��'�F�"��/E-��BH՚2��b�'�`< �h�	-��$��H�'H�u��'\M�B�=�ʑ�� ���d��'�5�a�ܨJ<p%���a6FE!�'���K`�f����Z'X8n��'�l�Q �ާ/�&)4Â�MVL3�'�nٲ�! �I�����g��Ua<8�'���W��t�FH�!OޥJ,���'��\+Ũ�e6 ���.<��!�'j��B���=,� 9���A����'_4��D�=lA�XvO�>��r
�'ώ���B:4ub� %�#�:�:
�'W��� }�n��T�@(� t�	�'h���2b.a��80e�ڔ2P\��'}��F$�M�������	(�0�'*N�h4���21Tx@���kC:�y�'Hl1B��H+�<���N�7g����'m�pP6
2+؉��@�+/|��
�'��m3R��(+I�u���ى%I&�	�'M܃����=gX��Ug�%��Ҿ�yB�X�`z�ȉS��
O�0S!a��y2 �!%�����F�<�p��Z�yr#R(
���C�IR�C��i$NA��y���X4��@�fW�<�4P�C��y�+�W�� ڕ�V�GЮt�SJ�y��Q�e��u$ �8S�՛��צ�y�D�F$��.�ҘFNמ�y
� �أ%�ؓ,(�%S��	U"O��!AIKH��☹6��bW"O(�!��Z
 *M9�@C�{�2���"O��5&Q�\f4�Q`�F��"O���`�S�6"6�P��87��axw"O���W̗�/�´{�D[�mѮ���"O��)�D��U�2�@���Xe�Ȩ"OR�(%f�5t��a ��'W+)�I�<٧��&xK�L���%_���#�J�<9wnI$RXh�ڰB@m��aFI�<!���9x�p!�I�Ь����A�<�2�� k��P�fER�@H���|�<��A�� ��!`w'�A����^�<P��& �p ���[( ×��A�<���N� a#�]�^F̑���|�<	��ZS�D�98f�ڔ�Ix�<��R�p���\�a�p�:�	K�<)�,��7�4�赏���@�#�|�<��#U�F�!2"שU�<�a��@�<ag՛@?(H���^���L�R��<�-��a�p������F {�<�����A����"Z�#�`� i]r�<i��C4R� �K�2*I�%��R�<a�	�.�<�@L/z~rA"�Y�<���Ϩ�&ܙŋP�cN�5����W�<a���)H�����)#��MI�<Q��m�Aˢ�$j�\��ΜG�<��a>uaX,��/]�2`�� �S_�<�u���b@ r.���bOq�<I����'u��[iIzB\#gdBr�<�$b�6Z�H�·̇�uQ��BuC�x�<�2m��}��5�p���IF���'(�K�<�P���څ��˄81��V-G�<q���/�nd��&�54�B���~�<	 ñT�]bS��\TpDI�b�<���G<ޅݶ �09�+J)#���ȓ8�^�0E��V�VP��V��
�ȓm`�%�ǭ�&)�]24'V�Ȍ�ȓĬQ���֡NM�B���z�ȓIo&���U1�&}�VD1^�x��CwĹ��-c���z+K�_�Ň�N�4d[T��iS��BA m� �ȓsO�tD� �����N�\��ȓ`;J�y���=^��,1'�ڜ�T��m���f�ΚQw��hUÖ"Tu����M���ɧ/�Hp�K�S�͆� T�YB[4�J��"�_$���t���!"�C�U��#4�C)����Q��ac�]�7���$̌�%��ȓR�䱐�1W�0��� `����a���� >A���g߇F�X(��D5x@tD �q�vͨ6�<:X��ȓl�iR��b!��5��� �4��L���s�*G<U��͚�k�N��X���40�/��	K~ :5$�84�ȓ#ma
G��/8���Bꌔ��U��
d���/�t��묈�ȓI�ް�`Q�@#Ѝ��c#.�����L��ȵh�4��	�t�K� R����α��K�+f!��
Q��<S�؄ȓh��HS�E9RUl�5�	V�h�ȓ�0|����&�1��nT��
e�������� �P ����@Td�ȓ\� ٫JGaH,�BD�;N�tM��S�? �츓�N�#\��CKP9c���"O��u�ٕ[��i;���M��A�F"O��p��$3`I��'�y�F��3"O��(b,�Ғa����F��5�B"Oҥ9�HT�cE�Xs%�F���"Oh�5,��?�,aB�&�
����U"O�#W�Q�M�T�� Ǧjw�D "O����,D&��m����	tq���"O5���
�B\`�,G.K��0��"O��#q�����t뚍���"O�p8��4�<10��&D5���"O�i�`m(H� �Ӊ�J&03"Ol���n��)$�,�0nM o�|d"Ol��2��$��0��)`���%"O����\t֌8�cؒt�B���"O80��� �z��7�<�^DjF"O��K7��p��k��e_��8�"O��
�C�-���ɖ�	0^�1��"O�@@`"X�/�2t�Qo��/Sl\��"O�,�VMO f��Y'��-Pl�1u"O�%!ck��0���(�X
$��u"O��bjP0�$�;NH�k�H��"O,9a��j� �q�֪E ��rC"O�w��r�&!���^�<�5"O��A)�)^$8���$�¸ڢ"O�ps��%F )��Y�Tl괩�"Oja9g��j����(w,fV��y���9�d�é@�&(`��?�y������2�`ڭ%�Ա;��M��y�gQ�8W��$4�(sǆ�y��&��b2H�++�b-"��G��y*�(k�0���!"���s'L��y2\�2�pE+���.w0�ڡ��.�y���,K%(�r�\�!�~��Ц]�y2Ybq��*�����Yp#��y�/e�~\F�+�nQ����y"�هt+�`h#	�.ˈ�q���y��پ�xϚ#�����̥�y�茄z3���&��@�ѫ;�yRC����+�G@�	�M��H��yR,��P��Y����I�4���Ĕ�y��	��Es�(ş���x!�Ѿ�y"[�v�&{�R}�	a����y�V#O��I��4�t�*�l=�y���1+�`�:�
I8<�T�#jä�y�Ζ=gX��Č./�,�jt�R �y���j��;Q-��"�jPaT���yN
�1ƴk��ץl�R��C��y2ba<�z2ˆ�dL`m�⋂�yr#�%q���E��Q��aOA��PyHU�C�Ɲ�A�*B앰��C�<������qIS/֣v~ ����G�<D��)I���CD�
'�L<�1\B�<	u�7t_z�+�%F=*�1ca�B�<)t�¹+�蒄L�@]
�Z��Iu�<���$E��f  �I�i�BJq�<�ծ�6$�ܡr�Z 9�Ƀ�]m�<)�ȃ'��c�lԜ0V��@�QR�<1�BڋE�0X�J�i	�̻]c�<�5E�;���B�`KFLJ�!���`�<�U�O"g4��G��.�z!�HZ�<�3��O����5	i�IJ�CO�<��V�x�8�Qϋ.1��X��M�<�$"C�j L����h�fP���@J�<� �M��F�um���G�#6��"O��
�K�$f "Ps���.��գp"O@9+F�;<&n��V��z��r"O������;7D�$B����A��P1"O�a�C�~��Y򌋥k\���"O����Ǳil&t�f.���6QY�"OR��b�)}�Pu`���6V;���"O�p�BS�F�n���l�0p6�} "O�@їD�*2�2�jT�9o�؛"O���0��=k�i eK�9,�@1�"O��I��=ft��S�P'(�P2�"OF�Baɉ4r`1TH�>@"O½b�	�7FF�0d��9��uE`�<!�j֖RMRh26�� �~�*1NE�<)�,�`�t\S.&R����<a ���t�
�fn��H�t�K�ga�<i�N���j�x�eQ3���Q�<a��D��u�R�G�!��8�ef�<�$ƀYM�,��#͝hbu`�O}�<	�l�:iDn8
GB�@e�p ��D�<���K�.aҐ!�" Yȣ��H�<1�IͲe���Cg���O���VOYL�<ISN�n���{� �C�������<1��R�<5�b�	�>����ÉK|}�i��DGy"Y6!�#:�<��L���=ɉy��J�ɄO4����dǝ:�yb"ԝN��ɠ#S���h���M:��''ў��IH��Փ��}�PA��(p�=�W"O�`F��@�i���[1mR��"O�	:�ƎT���⧤G�/R.�"O��޼+����4F;^��X"OzQ,�N/R5jU�֑QA\�;��'ўx8B͏�@��5S�*�AQ@�#&>D��z@�4@[:��Y�H[nu�;D��*���2ϸd��j20Y���9D�`SKA�q�T�Ɖ��s��Pq�5D���O�(
�&t��)W1R�8�d�5D�P1��=SMtuг*V/%�Du�u�1D����hld������lU[g�.D���� F.^l��s�8��%�-D���2a��4mJ�%�
����M.D�l��dǲDܺ-y��c�"7(+D��ʅ鋃8��rӏ��`��*D�ct���z����::���[K'D�رD�B�����C_Ga'&'D��r��!y�&�ӨB"&����	(D�t3(O��k���[�����$&D����C %!6��.�'�`Q8�@0D�t�i��_R.	�.ƸO�H��+D���$ǅ39�N b�ócc��9��5D�����+&���U�]�=�؋h3D���T%��@��7eWN���+D�7�]2<��iS���H���B6D�b�\9����F�O�D�(��)D��D
Q;Dא�	�ËL����)D��3�)K5gƈ�(�L����S&'D�\�d��?zf8K�H�~%�`�! $D�  �lTF<S"+E)wm�P��J$D�XZ�n�!K�2]�G�L��A�J#D��˷��7�� ��lLJ%[��3D�ās�K⬍�׌U�b}I�n2D���Ba�O�ΑHF�_�L`�:�1D����h\5,�h� T���H=A��1D���%�xҨ����5�`� c+D�� � ��'�
>��:��ЕR/�`E"O~�QrJ���h��̫1/����"O��ŋ�/Z[t�����f�B=�"O@��F�<f�NA[3�ݮ:{J��"O��@C�^lP0!#�H$&�dɢC"O��p O�~���)�=���"OXh#A�Sq�iE)V�Nv���"O�0�Wm\
P�X�JT�T� \�b"Ox-e�Z�M�2D ��F�~�i�'TtXIC�lJȄ��T'Z�z�'��A3����v�SIA�Th��#�'�&Щ�`�
��My���$G���x�'�<�	��FY
Pi5�� 5Z�`�'� 

UKR�!¡�Qh��
�'��e(� ��`�"�Qm�6$�	�'Ϭ��"\�U�j���ͺ/Sp��'GT�ㇱ:W�����X *�n	�'
�!��F���92��>�*�'���oZ(d���]�r0��'z��� e�f�
q�G�	5qX�'09�p�U,S��ZPl� F���'`����f��@WD�7&P�#f��'��;�jD� ��YY�F�\�����'J���F���찦�>CT�]a�'�R��cl**��1���S�>Y�p�'
>�I�f�<���+ �� 'L�[�'�摩�C���d�O'3E��'Un�ɗε��,��, 2l�`8
�'r"{�XPPJ�*I�
��	�'�H���")�F�#p�G-5B��1�'q<5�SF�5j䡐��:3��ep�'Ƭ��� 6 �Z���+�Zj�(	�'T0���-��09���ZCh�;�'����GR2m~��r9~�
�'U�Re���P�R�T�Ri�J	
�'��X�T�϶	G\]��N;f��a �'g���B�C��0�`�2��l��'2����-@�>���k@�:R��1�'4��7�ΓW�����J��r�'��Ygg�Y)��&��@ɒ)��'��uI��3�@�S枇0$�|	�'�ؕcE��H;X�8�w�J�s�'���a�'�"�$����<<u��[�'F� 	���DY�q�o�i�@��'��rW���q��ԁSM�U�J��
�'Fq�I�&S眱�ŢKb։�	�'l�,0���_��i�t�z��@��'hz�&�T�$q+C�q�n���'�>9 ��mز���B+h(����'�M��%ދ/s�Ȫ�'��\�� �'
�:C��>�\�t��*�r��
�'��I�C�P�	bD��'Xd�ȓ:��I[Bb�/�$�EÅ<[y���.�ą�2,��Tk|��^:2�ń�8P�����(�Ȅ(��G����ȓ֊!��Ă�rS��2��[|�Ҡ�ȓKXLEz%ßۆ��G-D.��e�ȓOP�Uڣ`��[,�mzc	�c�n��ȓ�.��w.D�#*�B�Q��|d�ȓ��xhDO���f@yK��H�NA�ȓ5�D{��=Il1�w!�=\�j��ȓ^�Abb%{b�)���<>�u��{ҹ���� HG�� �N5��ن�V��1��咂pѢuP`NŌ#��݇�S�? tm��G�N�:�$ Q�!w��ذ"O��1�a�!u���qh5lĈ�"O"�"#!̾k�T���A5�E�"O|}�6�ϐw)�1�4JA�8� �j�"O�酣 X!�	�	Q�Ƞ�"O�	�������6��uc��"OB;�ʅc+�H�T��k_��+�"O*E��:(T 21k��X�铡"O\�I���Ix�4H#`ɸ!,�"O|y+�#�S�{��;_$zQ�s"Oܨ�Q�A�.�X�jf�C�RHȴ"O@��"���j��a����q+��J�"O��Q��,�6�@��ܹ::P��"O��棏(Nm����Q� ��QKa"O"|���O �0�k�ʕ"l���&"Oj�"�!�?�=񨉯o��ţ'"O���b�W�Д���
��y �"O�dS3��w�����Q''ꌉS�"O"�)��)L-�8!�ӫGE���"O
	Q�BI��ܣ1+�m'�@RQ"O|�r�����Q�ىd�:V"OD�(��Y�T�R��&�-I�"ODEa1�*2�� b�V����"O�<�t�m�8[eo�-U��M�"O�X!GŰ;��E��'B�D�TS�"O�׍��<�!/N�/,By�'�?D�T�Po�X�b0@�A�P6�s��=D��+���T&I���ۚŕ��yr.J�X�� ��UZl�����y�J� F}H����5N�d��Ɏ�yRD�x�,�y��ș�.���y�����MXuO��o�ҽ9����y2��[���`GkCR�RD6��y��N%�.UR7L`����]��y"aEq��{�%�J�.%��F��y"dܨmV=��F*8�r/ĩ�y�B�(����,M�Iվ�+�J�y⮔��l�`Ӡ@D�Z��F���yB"�BBt��MZ;v�)uP��yBȂ�.�n�Ɇ�ݿ!Q�`�TAR��y���uY���IT#�������yhŖA���v��<�|��"���y�b� zҼ�a�+�����Q�
��y�G�?1���P3Tp+2�[��ߵ�y�N	�;�Ȇ�a� �c��Z>�y�@�'��Hx�"�B���e)��y��'v����@"޹@5J�yb�&cU�5*F@�$�������y�Ļ<��$��b�8?���O��yR��h&�9�VE_2<RE%�y�>aÒ@�%��6d" e���y�"�g�,�f����ĻBN�y�ɓ(6�&\�#бO�p;�ɔ�yb�!��Y�V�ȟ+l�z���y2'M�Wb�d˱�8Sb���7V��y2�մ6�)5�%"���K��y:<��!(t�9�T�&��(3E�$D�B�EX��L-�4`�T���"D��F�ʩ���I5�R�T�T� ( D��� ��nJJ��wρ=Uj�?D�P���]��\���A�2����>D����(ܺ)�V�@�
.L
��9D��yQ�0;��H�8�L� %8D� �S�%,ߞ@�k�;�(	@�E(D�� *���"M�|-�0��(�\��"O��ZA�\A$�)w����*2"OI����@l�!�a%�D��"O0�)�l	��A�U7(�)Ce"O���%g��,�&�H1�§��\c�"OJ��B�Un����M�<��`�1"O��e��\q��[�ꗏ	�0�"�"ON�h�Gʓ: b�#3j�r�y�B"O�X��'6>�\�C�)yəa$�y�Ύ�]��0�.Ķ=�&� 6���y"��4�uU!5�p�"䢁&�y��_��XZ�`��2Q���`X��y"��|?j�`��'��	��^�y�΅
��	��퉂�xAsl���y���~f�P[���. eS���y��J����I� Fi��@�
�y�E�2f��gK���<H���պ�yǘ)Hq�r�NZY�� ��y�I�>�Xq2W��w5 `C���y�b��H���"��q�}!��>�y2M�=~�: ��䊧j�2����֥�y�l�\ꬥ���ھ���g��yR�'�h�����
y���tJ�y�������Y�Pc�$iX�y��� ��p !�
AHc���yR�̪N���5+޶$J�L�I��y��:=j�)x1-�-#�`��� K��y�H�"8����E�+�^`�bOҡ�y�Ɨe�"Њ�������y�eH�dy D�b x���!�!��y�� *��A,��o �@`&C_�y����ǆL�[�B��e���y2O�;ZT�"�
E�#�
M��B�y"DB�hO���V	X8G�Lx�tH̺�y2���!B�R�`���/��y"�ۍL�l1C�/L�6�҅���+�yb֙a���2�e	`��&�Vȇ�~�╙���$)"��#��8y�ȓ=��9֡Ǻ��D�!�F(z�ЇȓG3��b�@���P������t�ȓ#Q-���á@;����h�8p��-�ȓA*��R�Ǉ)WU �����A{��ȓyJ}�T˽<�:��C]	��ȓ0��I�I	�R�tAB@��i|����L�N�:��/����*i��Єȓ^���PlY��Ls�P0*B�����z@���
=5?F�b�Ǳ;�d��z<��s����I �@��82�Z@�ȓo���Y%��7 B�u�U�S�P�:t�ȓo�� ����jZ���2��'~=��ȓQ�(��q�M�
	.�W��>@i�5�ȓ*��sv���h�@���˃GϼD����t��.ct*2��`t1�ȓ*��=���՝bE�`c ��� wx��ȓ{v"�k���Vኃ�A�7L(���䭲V#H0�xl��>,����{$��0���4f��=�v.#x�Z݅�VW�5�a-W%~
���A��eܠ%��B���ȗ%�h!��"ޛf���ȓt� �Q��qBL8�E��qs�܅ȓ#�(3f"³v��x�!�t(݅�e���А���ڰ�0�拷*X���ȓ%p��Vb�W�*�@�7C�$�ȓBj�UR%%N�|�����I|�M��S�? ��)P-p%�'��+�d�"O|M�ۉ@�|�%I�p�0�S�"O �A�-�"ʲ����S��@R"O�=ۗ���(�j���I�/�V��V"O���R*L� �s�O�Y�Z|�"O%H֤w�bd�'�m���"O��r��$������h�"O b��W+Y���	��Q�
��`ۡ"O�2�B\�_W�����"��2�"O6$�� 11�����.c�4�9�"OHm��,ڎ4h��s�E�# ���S"O �8w��+&�����Q�"O���B�!�F�#S�	��l�2"O�����T�@�F J��ü)��u#�"O��s��&�~ub�c	k��TxG"O\컐	*V"t����06��&"O�}��,+2w�m�1�N�Y�"O�*cTQ���ֆ�&�$(Q"O^�b�R���E0�g�P�l�"O���gVEr�5�u�L0.iXUS�"OV������6��F�R:t�4�p"Ox�P3A�.G��$�&��lJf"O�Y@���<"ܚ��;:�e��"O"h8��J�S�A�둫�
TW"ONz��4p���p�Ȏ&��ջ�"O���'�C9ݬ�
e2u4���"O��it��I��a���&�A��"OL,Z��e/8(!eO	����"On��BlQN�[q��#S��  �"O�GEX�q9�ɢ1dDIV"OFɚ'��%*�ɚQ�"]44 �"O:h�ׇ��0�"<��Q�.�T�"Ot,k�U<t9�`;��%Ε��"O �#������h9�B=b'Tp��"OB=�a��,]�z��+ҴKtzr"O��k)��H`�Y��G�L��X�"O\hd\�a�@��i�4 �D�1"O��`�-1�6t¢�8k;����"O΁`ֽׅC>�pAL�f6�`p6"O����!��]�ċ�B� ��U"OfY�p)gq�7�ˮ\zlcS"O�|��A��}�����3Ty�"O���CS�[!~ �`^�;1��sE"O��!���0͢ѥ	1 �=p�"O<��&
P[Lj5$�G�ny�"O��I#$�1d�}1�cJ�\�J%+��)���OD�T%� ��ü�f���ÝG�(�A�.D�x��˙�'8�h�C�' �hx��-D�4�&� �~tH���ߊP��5D��*�EV�Z����� Q�cj2D���IU�2�����.p10�
1D�tp��*7l1�0�Ȼ5���Ձ.D�V�K��A«�HJ�#eƭ�y#��y��Ĉ
5��7f���y��8��dY��2s�F����yR�L��M(B��(,ވ�g��y@X$�F�9AL0�o�2�yZ8Y��ҫO@�� /��S�Hi�'g�ѸOҿ�~�*V�P��]��'qf(��n�(��,!v��d꤉�5��x2�V*��|ؖ�ZKX1�DB��y2�
>�L��W/��K�ک�ᬘ�y�CK�-��,XcѴL���@�X�yRӾ]����Ä|�컃���y
� �3BeVe�8����_j�au"O\�:B%_�ݸV��b<��"OܻG�H�g��$��ET������O��L&�c�#��+�Xa�#ʍ}�¸�bk6D� B�jE�6�F��H�f�j�q�#9D�8"a+R�s�F�!Æ��`�9D�D�#��DE����8�ݓe�7D� C��} �*�e�4�C#D�L(cB��	$r��`� 搠�u-D�`a5W,�vtۧDN�O���p�,D��	0� ;�`s�M��TpQ�`/D���f��$-�IS6�M�t�`��$.D��8�LT%�������+D��y��M�$�@10C��3�(��(D�8K���A=X�q��@���bT�(D��P'ǂ4�<��ae:BfD��'D������OK$��'��TK>L)�m/D�xQ��þ`-"]Rf�ۋv�K��,D���"H�Ba�i%#Z�[FJ��b*D��@6˚&`N��l�ioN��qh"D��i���=�Y���ٖ���s��!D��ѥ� ���j�؇3e�����?D�97���і%Bq�		��+&A;D����ՑX��3RA�[ys;D�`R����aSFa�5K��Pq��8D�ta�N� ڬ� t�@�g��9�ы6D�����7&���1��5~X!S�L2D����������|AF���,,D����%? !5#^��E�E�(D� ���_/F�f�aA��'$D���ဂ*[�@�"�]C�-D�Xj�W�*ւ�0��HIAn*D�\qD�T�+�}R�%�2H���CR�$D��x����)/�-�0DA�w��釅=D�SPK#{ߠ�B%䞌&T�M��J6D��K�^4 �bm=������2D� C�U�n�83��Ě3��r2
0D������x#$D ;�n9�`,D�<Y��E<P�x�����+H�i`G�(�OF�O��aj^��`�U��0e�~(q!"O*��W�'��|2�-(�B�2�"O�����I+7����Y0���"O�m�d��>?�Ұ��ar�!��"O��Y�aD�0�Ȑ�C�� f��"O.xI�n���� N)M<��"O�0d�� ;�q� /]S1[P"O��ٴ��1=�l��$�e��qmA��y�p�l��E�j�:���K	�y"+Em6 $�0��h��٢��V��y�u�Y�@�=g�|L@���y"�2%�@�Ä�_��5��l���y����pdn�9%��D0�f����'�R�'�B8`��*,��JP˙����A����OΣ*@��#9 t��?HlL#�"��<W��l�j��E���%3I�O�<I�+J�%^X��o��pu��b�AQL�<���ϗ:0T<�s�j,�DG�J�<9���)�Ā��d�D�>*�]I�<�a�$��I���͋$�pu�3
VH�<���L��yy�e������D�<��+˱7@N�#�C&5e>���g�i�<�0nړL�nb�Ģ\���T��d�<i4���2�8�5"��0�&X���Gb�<�Q�A��qRC�\83hpv��y�<� ���uc�.��Pf)"�2�j"OD�*���_>���$�Hϔhz��d�O��?���<OV��k�!��A٥e���ȓ����C�4,�I��	6��ȓx�R���WHĔʥn��]B؅�B�"8"���L��[G��R<�ȅ�f�T0At�\?<��1Z�ޙsHH@��Z�8ET�k��4S^�քDxB�)2��8 �	MQ�����G�<��.I'uj��zCi��/a�	��nWC�<ђ�<t,m����8qFՠ�K~�<���
*Q�`��2y)�;oXt�<i5��f�:m�ï0:ppY�Umn�<�	�
zB����*@(f�д�Nm�<acǑ�a��q���S�H�Ppp$A�h�'z�Ik�������@�&uz�	�Q?Ih�ȓo:0aCIѫ��p4���Q��`��	B��ȟ��Q�vE#��J&C����8D�@���t�$�� �:t�nys��7D��T��>vǼ��� ʴPMT9�7�;D�H+AH��
S��T;����a$D�D�C�Y�6��%�
} GC%D��Z%CB�R�lrwA�V�"0��$D�Dxw`D U襤z��O�"a�[�(#D��1�j�C�l�k���#{�
p��M<D�8� "Ҟ"b�0woO�]�,����-D��J&@�3b����P*R�L�y���(D��Y�o��^��m�s�* ����(D��� \"X␘21`�gqp!k��%��蟆Q��dߠU����%)�Uj���"O�����W�y�
��VN�\���a6"O�<	�'�l����Mt��p"O��ȥl��]�D�JԢ�
<���� "O�Q���M7t�~A����&c����"ObUp��2`�@�P�Z�A�<�ʒ"O�l��B�u�!��"`��T"O��:�.�B��E�D[�h�"Op��g�6Yd$9R��$`��"OX�11�0lo�A`b؝E��"OjɉsD�e�.�I�
A�HXQ%"O���Yj����J����n��y��W�a�Pt�1`�qo֤�y�$�E�0#5���(���(�x2�'�"��!Nf����J�	�f��
�'64��$L}ѐZ�c�pvP	�'��ӂB�rz~�+�x>(�
�'��H��C�<brH ��
H?%��	2	�'��Y�w�^��[B�œXX���'��H$)�5��0��$�=g�8�#�'�����c^�8�hIR�&��,� ���'�h��j���$qCD	�<��	�'��؊U��=1*%��+OJ�4��	�'�"�����8pLq3�ˀ;=��	�'�� �r��&U_�����2c����'��*)Ƽ\��L
"G�v��'�Te��m�~Sp(�g@�k��
�'`ĈVg��*-���X��p�'f���Ńw²iscI�M�^\��'لPJ�L߈�:��잋r�����'��A�u�
�fzz��e��3�����'�t,)&n5~�f�#$.Y8%.> �'Z���i�XLh2� jX��'(�@DS�|��� �&D�	�D٪�'<՛�⑚H9:����R�i�tQ��� ��%�فk���ۣu�2�"O|�Y�e{�
$�OڎV��p3�"O���B�o�d�@�v�D+�"OJq�R�#m��;4���,�\٧"O�9�̗��X� &K+j�fY�"O\���S�L�r����v���s�"Odh�"�d��5R�
��}��"O�9cD���v�pe)䌇u0���"O�Pj�����}�',��cy�"O�-�U��!D�jd��MU�~e�"OT��6�ަGd�Q���T�"O��W
Ҥ�(�	cI/
C�@6"O�i``��	Y~T�¦A�G���a"Od�[�3*~
ɺ%��#�kO"��@%at-(P(��F�͂n��/H��3�O����@����-ω��@�"O���zfD5��F[抁�a"O�q�t�����;��&�0��"O��y�eæQbP35��n�8]�E"OTY!�;1��$(�Ŗ$Ct}�u"OD��
�P��d�*fXVh��"O2}�fGH�'�Z-�#+ig��ɔ�:4�4W.ݸN��X�1�O�M�^I�6D���PM
J��8�@O�=|��5D�Īf��%�B��2�"&M1��/D�x��!Z������O!,2]�à.D����G�,oh�h��)/j�Q�j-D�����~��0w��z%Z����v��y���O���S0-�𡰓M��4:��A	Q2O�!�DT�i8�ܩ�鑱P���I�!2�!��n �zìέ+g�ȹծ;Bz!�$�n�.T�Q��;r��I��mJ6X�!��
�#AL��t!�'(=�U�r��!���K����	W;CWfy�S�I
�!�d�{�z����aF�I[`�=� ˓�?����?�|�.����8@[zX	7�Ԁ7,M(�A��!�dC9u��-�q	�3'��{& J	�!�ߨsT2m#Ӫߘ�6�f��b�!��9z��� ��rԴ�"�K��v�!�D��c���J�e��@�r��XW!�Ϊ�4�B��0O$��G�@�X+!��D$H$X�*[��-�ӥҮC�>��?1���?�|2/��$ �<��QΑ�&���%n!��ރN�L@
 �Ϧ=N��!���,S!��"�X	pRn0'|Kp��UB!���%tj<1eC�`!� A� T�!�X����R�T��u���8!��W&\����wt�)tO��_�!�D:~2� a��g�˄CO�S�,�O��S�g̓D�8��ɕ�tV�ѪD@R�N�j��ȓd����l��kM
	��gX(��%��0Am#r���RG�K��m��uCԨD �#����׎���L�$Z"#Cv��r���$�ȓp�z� ����Jޕq���.�`�ȓ	Nt��#�ˤj��aQ`��&H��`��'<h�p	R�km�ŋ�@����ȓZU�	&� :EYBe$o����ȓ6~}0ceZ���%���g�8�ȓy3 @c�ʓ_a�� 3-è~u����T�iiǈ�.w�d�e@X#"����ȓmyf]�p��N�Z�&��`D��ȓ�dz�ɇBhԵ9c��ȅ���?�6k��r�
��HԢh
��C2�W�<� �T�4'�0"��zt(B"�*�e"OB9:po62����A�W"5|:Ԙ"OZ��`Ǔ&Q�J�s1쓍kt�B5"Of�9�W\N�P"J�1]荳4"OzM�`�9�:����oZ��1"O�U��W�<z
e��g�/(u��5"O�����+>L����C ><H9"O|X���o�rw�_8_����"O�LK��6 �>%XCE	�OGH�2w"O�	yE��;W��4u���t8����"OZ�(A��G:�<)��_�{"�!��"O����"!>�x�惷9�J���"OT�(��C0T&���v�SB�']ў��Dk��Aj�`���3�px�� D�4�O/G�ޥ[��%H���E�#D�H�TF�>hR��D�<�n���"D���v	��S�̐�Ѩ|�FaS� 6D��㐀}�r0s�H��j���i��4D��q��P�>�X�H�l�V�`o1D� 3�&J'Q��%�dŎ�T6�uB,��� �S�g'Vz�у8��Ī��а\��C�I�_:�aҚcX���"�$9#�B䉦?x�I��9]��k��2`��C�	(9�>(��/%l���é&a>C�I�VP� ��( ����%F��z"Oz�Q���\�{�'�%*2YKE"O�@A)�(�IeA�#Rz�!���D0�S�dO�	�H�#���rS�-3����y���%���;��Qrl�x����yREבNw��sE�<݊�ʡ�Ҽ�y��L�9��-҄�Q�2� ԑF݂�y� �<K��s��`p��uF��y�bQ�8����nY@��4Þ�y��J�d�P�
W�6�J�kGJV3�y�h��0 \�c`C��E�%�V�ś�yҪ�F$f}�S���0O�􀱋Z"�y��^=6]|5�7听3BX�ˀaQ4�y���@�Z�A'K� E���"�y�&Ĕ~0�)�i�9|?�H۷GP��y�Z�*�a��ȏ|������2�y��]�X4�@0�1+�|y����y�N��
�C5�R�5�lA���1�y�&B2���͒�e�������*�y��#��)��C�p���O� �y�*D�	¤A<-0Iw.N(�y�K�
f�x@7B�,JVb��B�#�y�㕡l�¥I�� Z,8�X�yB�ܒ`_P0�c��(K�8��`��y�.\�u�Ъ�!�o��lHwL��y��ϜNv���VM�|ޕqAE�y���"al!3��7�.!fG�>�y"�5|��)�ǍU>z)f�@�y�V�/}���l�WD�Q{�����y�T����'��Q��UC�4�y��<��c ��S�,�Ȇ��y"�1���#���-���Ч+\��y2��)/���
ސ�C���y�(� |�X��G��}n�P����y"�t�dm���[#zl���sfV��y�℩TI��SO�#u�N(�eZ��y��O����p�-���Py�i�2>�v�� ��T� Ӕ�Cl�<1�f.H=B��`��}�5��Bk�<�4*�InTi��"0;���T�M�<� P˕	��7QZ504@�0�Jx�"O����Ӕ�z��UI�3` ��"O2�"e��m����`-�7���b"Od����H2cY�t[��lX�Y"O:��D���P�xVHUS�"O����ޒ\� �J3C:URvX8�"OF\�&O�<t�0 GY=ISމ0 "O��C4COڥcF�ܨ9N�M;�"O>�h�$[lpSb�64�q� "OTP�"�Q(�pp$�]�V�j2"O���I)|���[���$s�L���"O����O�&1٘�A%#�#ȨC"O��S̨q�N��bL�n�)�"OF�j6�VҸ ���9:�<5A�"OȜڂ��]�t����z���y�<�3��!J�2����5ol��To�P�<a2+U�HH�����}^�P���O�<�Ӡބ�� r+A%�&�9�-g�<��/s !�)�{�xxB��y�<�3��{���+��.�X���$s�<��(\�%�ؔ�B�֭p̔%�Jm�<1@+)=��ЬVM��x�AMj�<a�'ƻ����dO?S�&(�DnTo�<�횉yp �@p
O�6��a���G�<��Ή9n)�P���5@�0�K6)�Y�<��m�3
snxi��,(M8\�V�<郡�5b�ѣ�$˩|Ոa`E�Uz�<$�Z�(��B!"h��1��y�<�r���#+�Q�(ya��Y�<ᑥ�:�x094��X�(I�E{�<	��B�n�h�.� �dD�Q�w�<q�߫A����	D����I�<q�!@, ��b%B��Ӛ�At��Z�<�e"G)t_,�3�I�� 0ԃ�p�<�V�ÀZx`-�ƁM�"�����Om�<�E�/@%b��87����&V�<!#`�/JN5�u"�-5|�pb�(|�<A2bԋf�$C3G]�86�hR�M�|�<��HD�rUJܤ-?��##!�dܒ��a�?qty��d%C�ɲ�b�;��R��Ѕl��}��C�ɯ�A	ѣ��8������(��C�ɢ �x���
oց�"��vC�ɾNL�ej��WSx�Y�U�}&xC�I��ɱvh��`y��Af#���*B�	&*zx��a)ˌ}�  :C�	�>��k��S1�43-�?0�^C��ƌ�2bƓy�t���A-v��B�	;������&5v�t�w�3k¶B��}?�Ep�Ɲ? (>pW�_2�XC�	�n�J��b�Ԣ���5�
�8�PC�ɆG�l%ჃR�q�
TRf�:�>C�4S��#A��D��� p`ڑq��C�	#6B�re�R7����!·+C�Is��e�퉓F���d��C�I-=[r���n3X�΄���ܘv�JC䉑�
�@��< :��0��b6C�I��t� ��
im@	���Z<KlC�I�>��Qa�}
�KW�ZO��B�I�/�Z�*%cǈg1���Ǚ�>�B�Is�~l:���\��t����?��B䉯S�3&�Rf�R�1#T y����;ĺ*6�U.����K$�!�$ːc�Fp��^g�:V�F�`���� F Jg ���(��!C�#|��"O�ݙ�Mܦb��@��ΰ:2U�C"O��8��һ~�er�j�$,��4��"O(h���O@ 隌1���#W"O =�E��{^�Ź�!�Y20m��"O�@6:�N�����?"AZ�"Oz!b���'p/b������`�a�"O�\�&�Ab9�d)YS�z "OZx���
T�}���ǜ4�v� U"O�
%�,�c�"�Yt"OR�)%&�r�J���'�2�z�"O���f	(x>��g#~�C#"O�����;�8f�K6X����"O~�ZCʖWkzP���|!C!_�X�!��:&Ҵ�s�Յ`��4�#�$D�!�d7����[�H��RK�,2M!򤌳ET�8�J��G]~ ��)�y�!�䛤N���@�K�m�v����\�=�!�dB�����F�>p���q&�+�!��I#:Z�T�-6%V~��B.,FU!�$G�#�(hQS�
h7=�� b!�D��a�� ��c!�Pz���%I�!�D��+����#�0�� ��&D�!�d��~�����!J��X �T�q�!��:��a�P^�?���1d�v�!�Gu_6���F�,�s��>!�D��`������x�9��щ�!�O	:��HY�n��tyT�f.�E�!�S�Q������	not�c�J 6�!�d�7�h�+���pf���T�$�!�S�߶Q�rm�2GaHč�`�!��B b�#u�� abO�N�!��	�f ��j.0�:���$�16J!�dM.g�ě4��ߤt¤�3GF!�$�h���ąl�b�a@2[�!���"t��	˰W�	Yr �a�!�d��" ���!�=Lj,�# ܼ�!��i9��2�8p���0F�!�ǇTw�����L�.r�r ��Z�!���=T���Po�7��!��OG �!�䙾|O��z�a�><q��'�@+go!�$�M$���/}��̛��V3Z!�TLdbT��-K�e�D���J�:/q!���Z���c�d�"B���ì��8!��%��Æ����0j���(!�DΚ]K*�I� -������+'�!��ڞh�����B�YrE�6�!a}!��:\U�!" 4eOn�����T>!��c�(�D�Y/�TA�!㔚P-!�d�&��i�l��n���t��!�$H�'G8��%�/7�4x�@�5�!�V% ��h���L�J8QU��!�!�ę�X�V��v�"� R��6Xq!��d6�-t��n�� �0"Ox�g�J�\^�ջ��$F�z<�1"O.P%J�r�lh��� �>({�"O�Պ�Jް���w)�V��	X0"O^�(S��yZ��7ʟ889��"O�9���c�̼�V� #+tQ0s"O�A��˓�n�A�I��d��+b"Oơ��� 9a�x���M�ih�}��"O�Q���A6C�0U��� uW��r�"OR� M_d8�$�E���"O"E�#��0]XZ<��ό,\��b"O� ����R���pT	��Dx:h�C"Ol�f�2`ڌ)�J��@�"O��M���Ks�s���m�<Qt/�6�������>x�����i�<��L��
��Do|�;��
c�<y*ǚ6kl�3��[	9�	���.D��YB�� �T,�"b���}Iw'9D�Р�&@5�,�6��O�����$7D� F�*ʬq0�7r���A�#:D��P��Kŀ\��!;2ry��7D�,b�,2Hb�5B�&ޚ5zL1�� D�8��Gm��8!ǗB��!��=D����K
&�-�wΘ� ���Q�a=D��Av/�/�����B�S�R��:D�\�A-J�g��J��@�ź| ��9D�p�CK�8eN�Xf� (����4D�,,}��L"4��5��d��(��s5!�d�
�~���;JI��bs��_!�$k�1ȗ'E��GFP�o
 ��"O������sx�D��D3l�g"O
 ��'�-rH���-X�|�D܃2"O�9��CV�s*`�ѧ/o�&��0"O��u�2�*��a��0!c�!�"O~sҪ֒)�@Pa�>>P��@�"O����'�<J ��Q��<+j���"O���TkX�M�F�Cơ�Ex���"Ox�"vl� $L��i���w"O�����orޱ�"Ύ�>a4��6"O����1dd(uH�;!B.��#"Op:P�WJ�X`B���v*�a �"Ol���%ػd����:%32���"O<4�mT(����������"O%Y4M˸~��9�c�؃h���"O\��𥑴��qJ��VB�D*5"O��
 bŖTP��>a�8-�D"OND�Q�E$e�rY����j�"Q"O:l�F'�Q>�����'���"O�h`��� �����B�	Ǆ#5"O��q��ːSj�Q�f-��Ț%"O֠�`�j 80/�3��U9�"O6MЂ��5C�(5�hM�M�ad"O�@	�I�F,��U�	}�Ht��"O�]��+�< �}� CW��vp�"O2�K��K%�r������tRu"O$1ò�Z���|�t�G� =$�"O��BB��f��j�7(����"O>	�D́8�x������	B�"O:U���_�W��U��*�0v��"OI
䭟�0���AK̴N1ΐi�"O�<j���-58M���Br~壥"O�����($N�C�F֐	�,��"O�I���W�\� -���O��ִ�"O(�҂�ߖ"p1E�� _�D p�"O�ɀ'.W .Ej ��bD ^���Ȕ"O�1�l��bӗ�Ի�,�s�"O 8#tሣ_p�`� �O7J8��"O\T�c�Uxθ�2g@ۊz�}Ku"O���TM�Y3����x^�X�"O�EV���{�H�ԯ�uan��B"O�`2T�;O0���H&M ��"O���Q�]�w露��ÿ+� ��@"O��2�K7s�2|�҄ˠL�v@1�"O�@WJ׮<8Y� .�޹�"O �Ct����Z� L�h�����"O� }���:��a��4�4j�"O���S�͢7K��U�ä.�T%!"OF��&��2u�EQv,�b\
-1�"On�����X1q�/DlQ4"O̰��K�Oc���b��e�w"O����9,#	�t�xղu��"O�]x$G�'"��̑�� 8u�""OvP@��>wy�$!"	����t��"O����Y�2�.	��<0�!��O�#Y�iDظ3��5��N��N!�$�i���G�W*�� G�Cg!�DD�^��e8�a���ш��kV!�ҵ8
�ó�����X(����L�!�d�n�I� O+�u���B0�!�U�9�JL[��;Y� 9��C3�!��k��!Ȯt��`���A�!�$�R�m鑮�9y�i�2�E!��`50�I7��zw��8��[:�!���id���� c��Ǵ�!�d�=8*�x��ߘ`[z) (�/"%!��� �����NτG�h�	�l�!��t�L
�0,'�Bv%�x�!�D��B��l�q��ّ�+�!�D[=K�.-�ߣj�p����;!��F�3G�� e�\M`3O��#k!���L���$�/o?�lP��I�i!�ӄUJm�礉�����q!�$֕�½y��W;"��(B+EW�!�$�s;�AڳC�)�}y��.�!�W�z�T-�D�X"R|#F��>�!�d�C,�%��I�k@,��eJ&~S!�D(Baެ{#Fܧy���dG�fC!�$mX�;"���qcP8���]�q�!�d���`Q���+^���C��>�!�d	Ҙ�7d�4�{fA6Hۡ�֫ALy�fE��XF4-�an��yrk�#j��3oЕIJ�L8`Hċ�yBgM�t���W�GB��P��R�y�뀸D.���2�95�VqPt�_
�y2��;�nd�ĉo�q�SF�8�yNW��4�A"�w�i�BJ���y��D(�nx��=M8A�֕�y�P�^��;��.Fh�c��ȕ�yҌĒ"�J�b�DC�(S����L��yb$��-�����Te@qQ�^��y�B_�#��O7 x0�dɝ�y�%_|(�D�̜�=�*M���F��y
ǍY��N����ȭT�&	�"O����Ȝ�N1�W�Y�9�fȠ"Op8�1ER�R�0hi�bPfq�aB�"O���E�kq�5 �	uQ�mp�"O,�Å&�� ��C�T�[KP��q"O���ACU8X��Zt��)
>d�XU"O�@A��G�FJ�qkg��o4�Z2"Of�p�$X�oN4hb�:&�(0�"O�	�NZ�n}$LI6�����R�"O�P��`*Hz���g�� ��PW"O��r+�Cs��C
S�nc����"Ol��䤇�dڶѠԉ�6 T4<H7"O��B�$O[i�4c(��0<���"O��E�#mB��橃�����"O* ���	7���q���8?f�<9f"O�E�
�%&RZ��hБC�b�8s"O��څĖ�m�6����ѧI��I��"O� 
D���G�N�[�,�T̲��"OF�(6N�#-�
��KI�=���Q"O��R�/��"ky�*S�@�騁"O�ԈW�ES©����1�޴À"O��F��$B��L�)E�&�J=�C"O�̳sA�@�X��#���6"OXy����K�`Չ�6[.UX�"O��ka�_����g	�
&n�1��"O4[���0�QE隚k��P"O�\�c��$��iwf�&b`�s�"O8$�e*�p�B���IiΤ�1"Oz���6TA��:Ba�OI*q"O� �bU�<�×���nd6��Q"O���M�r�~�� V-�<�0"O���`k�  ?��B�a
�{Q�� "O���0G��f�:��+;�T�e"O�Y�f9=k�D �B�)�,�0g"O����ʱ\p�1D!C;/!p��"Od��O�u�� ��S$I��a�"O��{�N�em$i�����Az"OY+�蕥V4�=S��D!3���d"O>Z�ǐ7X��B�@E�K��x�"O|��')��A[bizD��X��I�"O��v%Q8S4pec"l2����"OZ��T���&Bt����S��\Qd"O4��`b��*g��C7$3�"p��"OR��p H�_ʄ��i�-P�ȜRS"OjY� ũ0���H *=����c"O����Hل
T�詓�Pk���AT"O�)u�[UT)�Q�F�<�Ɖ��"Oꌛ�#A�y��=Є#1B�x�S3"O�iɃn��m�<H#�Y;v��I#"OPI��%�� ���F��d����4"OD��W�ٍP��%+���8��QY�"O~�x��^�^���g56�@�SQ"Ol�+
�.��p;�f_+t���c�"O�����p��5D��!\��"O��k+ 0?�͛����vJ��r"O(y�f�WiA��х�?",*�� "O���Q��� B�(�`��"O�EC�d8�"p��J�v$�P�c"O���׎ʰ!&Pc`�֮P7��i�"O<�Z��'\bP,I���N��T��"O���Te:�vEK�S�pՒ�"O`u`�L0e"��D�-1�R���"O����@	Q���3�%��$�B�H�"O�i�b �������x��X
�"OLz��ތ;L�5�B [xLy�"O �*�l]���*�'
qN4�"O�`ѕ� 8�����Dq�4�v"O�<�a�~��p��ʈr�����"OL� �ߥ:�|$@DI�a�2 B"O���"��#]�lq�(O�@<��8"O`}P7�Y�8:"��A(�w
x�r�"O6��!2L����M����ii�"OF���L�F���;C��4>X�@"O��
�w���Yw�ŢO&0U�"O�������kv���
�Xʓ"OP�z"��2vpx���[<~ VM��"O Y�E܀$�e�����P�$Q�"OH�Pܑ|�ra�<�z91d"O�CBi�u��S�Z�����"O���A��K�t���^�=�~� �"Ofub��U<hx�G�`�p�"O� �L"�J 9{�|!F@�l:�ڶ"O��H c�$E)Sƀ�&\��1�"O������;龄�&�O�|�"O�A2�e1Ob��0��R��0A�"O�5�����4�pC���c�>誡"O��(C��-:'*�I e��o教�"O�S��D�<��ؑJ�K���K�"O��B���"�L#
P))C�+W"Ob�fF���<xI���j0�հ�"O�xK��
R�Eg)��%r��P"O䐊%O@�j�Н�&(EN�飓"OBA���&D8F5�D�Ⱦz <Y�e"OF Tg�f��,��'��x1�"O"�	4��?J�6t��ܺ�|�	�"O@ic��/R/,��E�gT0���"O�|c�� ��e�u�]�|;zP0"O�aсÀ�~<3Aځ2HD3"O<ͣ�+��*.�A�B()��z"O�#��"'��)"'�[�>(: 9�����OO�q����E.O��P��9���a�`\2��M
�#��ZtĆȓ!�r�(u���*.��Ʀ�$~�ұ�ȓ#�$��ǜqV���$�^�@��ȓmo:��G
�%��T�#���p�M�ȓZ��!��/�#n�Zi�G�������ȓx�ZQ�7k�?W�$qtc���ȓ�� 3�R)$`̅A҇��5㪜��`�t�$b�y)�$fԆȓ	�ÏP-���pC�EZHn��ȓ1�����K<v�Ј�J�Ma���i[�T��(;��,�H�=I�6E��X2�����X�O��#PK�1/��	�ȓl��|�7���t=�\S6H��9#R��ȓ	��P�DS� ��1�*ƶԅ�4G�<G�o���  1S���ȓl*��)&:��ͱ�gN�q&��ȓX��(@���a���$LS(k�\�ȓU3�T���KݤxY'�	W.��ȓ}1�Q8օ�o��Q�*��6Ͼ����!�g��o�z0	�%�#ǖ���8��	��-�k��	���ٜO��Y�ȓ:ӄm�Sf�%U�"A�k¤5<A�����H��V\N�t�W�D���soz�(�G�:5�&m�o�X��d-�4r�@
?>tԘ*&�C�t~(�ȓ5YB��A�ؒr����^1�v��|�aj�-K� �_�J��ȓUOl�X�׈�x�E��a����CyTسҬT*]�F��!:%�ȓAI�QcT�b��	���1�ȓV�R�2��A�1NƹY�)�;�؆�Fh���h��.����m��e
�����Ƶ1A�Z	����nZ�L����ȓn4�i�va޺R6Ќ �	�6��܄ȓm�jA�8sL:�����a20���[�h�b)>T�[���5w�Є�LۆpSB؟"
{M�g*)"!���F�=�t��������"!�ܫv�H���	c��ipK\#4#!�䑺d D�� �JH�ErJ�i!���;��K�,@�|P �c�Kd!�d�6"k�*���`�J8H�:%!�95e: "��?�&!�w(؎U�!�dY�f]8C��L�[�Q��a�$m�!�� ������%��dD&"����`"O2��e'��tYPPd��$3R"O|�!,�?^�� ���,j�f�#�"O���§�^�`Vb�a�ൺ�"Oy���Y�8�>�����7���"O���ekǡ-�r;t̋��T٤"O�p�/�-x>6��1m޺˖!R"O��YU�րPDHREF�6r���R"O�T���� Ǡ�����;]�DMA�"O ٔ�\	pL��ǭ�2�.�1�"Op���ҷ,`�ta��"�ZPQ4"Oĕ��-G	/�� ����b��Q"O��P��B�:�(�DT�GlL`t"ON�� �^_N8,A-�#\�\1`�"O�1W�μ@�L��7ܰ�|��p"O+%*�)��[:0t��2�Am�<!�k�%]�䩧-�w|�A��l�<yp�D&0Y���T�&m��A��B�<ARKY�^8VЩ��\�Zp���%e�h�<Y6#:[F�9�ը~��`;@,�J�<i�J]�r��J� '!	�c��M�<!��2n�̈B�E�)� i�0�Q�<�����x�df[8�ڤ��k�q�<�S`�)U�����^:�2m�v'�p�<�&AV�w�0��m��Y��i�<�#�z��!�����y`n�P�<���~]�D)�%���T���D
J�<Y凟2��C�L��X�I^L�<��Fp���Rv�+�Z��P��E�<��$P��yf�',:j-��Hf�<9��6ZA�mŨX-;�ٓ��c�<��X4^��T3T�Ս=�����^�<i��ݲ8E
S�Ř�>����u�	d�<I��(F����(ʛY��d"�c�<i�
��,� �گ=;�%�0n�Y�<���=p��<ej�}����D��Q<���C�����Q��Z��N�:��q�ȓn�}r���Y����Dȑ&XZ�����?���	 ���ڑ�S�`�*!�'�}�<���_�\��q�E	�K�AuC�u�<ѳc#{�$�8�ُAŶ �v�s�<�b��Rc���h�N�$a2��C?��~��y"b�T`�h�%RX���r�<�y2��~P��G\�0�׀Q7����HO�c��bl[�An$��:	(X�S�<LOT	z.O���o�@]'��fD8j5#
Pb7m��Aa�'M؁#c��g�PZqo&!���������^��C���M���D�4[�!�$ GZ$I���҂.�2,�&@8�V�@E{���0 �Q�� ٵQ!�ǃ_�g!��`�,!��a�=�t��cH2KI�B㉵
XFMb� D%kD��3կE9Y׈B�	͟�i�%\lR@� N�4�D,�t "D����lФi�!��"�	$|>�"�$?Q����������DE&�x��7\̀!y���yb-	� �H�Q!cƷAT8�pA��(ON��DE�4lȔ�D�r:p(c�ۆ3!�D�27V�=+"��Vy�"���:��@��F?�;F��D������mnB�	�:�xA��2��<����*�6m$��a#U>w�0Ԋud	5�Ν V�)\O���=���V첀�@"�v�|�� I
R�<@� x��ɳ� �n.S���X�'`�xb��,�:��jת
����Q��y
� 9��1˖	��j�<@$�G"Ov8���X=D���$�ԧm(��h�"O(`R� �Ѐs��ѝ7{q��"O>�cgE�}B<y�6����f���"Ox��Ԭˆ.lđ��nU�q82"OT\�G�,=R���f�Ȕ/�<Z"O��sFZ[ΐ8�fW�{�}�G"O��񃤄�{,,I����7:!��"O�#�,Y�+\�����\�S1"O:x��%׬�pk
hC"��5"O�ب��"z0��g넚8K�1Av"OT��E�1`4�d�V �.2fI"O0��H�4�8f	.&�1
e"Ot�"���uUV�i���	Dv,�"O�	���Ih�8�Sd�
8e�H�d"O�H�(H[t@���0VT���"O�<#�哓w�]+�DJ�I���b�<�T��E�<��1�z�H� ���D�<�p�&�����D��v'j� DK��<����)��a��ޑ\z��g�@a�<��Y(�`Isg�tB��X��B��/~w��H�-��&	�Xs I,0� B�ɷ ��ha�[yT�P���
#:�C�	'ZCz�Rb�\�C7��qREP�aZbC䉉$� *r�XBne`r'�$La�B�	�S\�8����@����~��B�I�3̜!M��<�T+e��, U�B�Ix��������ؘ䨒�W�lB�	�\BTe� .ό)M��K�8T�BB�I3	�~��5-8/U��yb�R�tdxB��~ҙks,̰'2��Bp푏C�	�W$��&@�=Pr�z@��{��C�	JeL4���*}\@���=R3pC�I�u���bPu���$`�^t&C�	1���M���ÓI'>C�I�A�q���&��6��HKC�	3~������R�����ŌJ��B�ɓ}���X�	( D�A#N&}��B�ɪM�<Q`Qʃ'@1�E�Q��"��*D�` a�˻}���+�$:��a2B8D�P"��\�&��T�](l���3D����ˆ�z�,Ě,�7�4�3�e'D����?#Y��
b�N�i
��%E)D�x`��p�ݹ�ˀ:�ؑ�a;D�T ��5(&�+ǏI�R�6I�C8D�p��ծ��0�E
r?P�8�f4D���cc�']nz� @D^��H����&D������S� �`�&$h�#@2D�x�	W56���L؛6�y�D�0D���7J�5A��$��&�W������-D�����;������Ȉ[�����H-D�HrԈ��s��g(�	7f���#6D��ْKEILP�%+�#.�,E���4D��[VAR�O4d�!ۀt����.4D��pF�./R�AS�T����W*'D�X�A%�R"��bF�Աu�8R�B#D��B�,-��ň� T3��m+�� D�(��_	lX�А�(҇��9�-1D���ME��IA�:X����:D�4��g��������b@92��,D�����2m���$�M�X&�Qeg&D��� ��7:�=0H�Z���Q�$D�@�2��gX�xBܗ\ d1�"D�0��o�&�6���٫��  .D�� *�P�{Ů8 �!O�\�r���"O�!�
I %��U�� @k�\�;�"O
���� �VZ�9�@�T�s�vD*0"OXI�gчt��1���z%�"O����N������/�Ry{�"O���� N�i�N)�؜g��e�"O��kT��*<�,�ir	�#{Li13"Od��U�\@���B.
�Ck0hK"O�m���_Gwt���W�JuS"O��+@�A�R�2ak^�8���RD"O��H��D0D�i�lϭ�x�Q"OZ}i��BU�$% �%|<1��"O��Cd�̣�i�>]PR�"O*��$lـ|��UrԂڦW1�ڀ"O���2*@�n�H��шN1�X`�"O��b��2z,�٫�^"�-�v"On��fNs�����j�-Ƽ�R"O��ܖ#s�.��c�!b�d�C"O^,#��˘�hm�Eo�!@۔���"O�q@�k^%w%�|��эb$vU1�"O�(�d�Ό#�.�D�t�R�"O��ʳ,�9ZZ2��-R#�@݉�"O��d�l��I��	�@�4��"O(qT+̻<��R�g���ʸv"O�D�q䎦 ��`���-(mpu�g"Of�cv�J�HW�0�gH�%�8XR�"O�`�
>��� �)psn`�#"OH����<e��Gһpl���"O � V/R5fL�JǦ��b�`�u"O8� ���(_'�Ars�M�lH�"O �t&�:jg�Ic���-�Z��"O��;�d	�&�i�g�Ikd�'"O0uRPJq�UkT���9�C�"O�\���"_VЈE$�ā�"O�x�\$XV�ɪ�M�Nm�)�$"O���'�[?���q��
QO�$(�"O��P��ם1"i�#�A;��� "O U0����l��@�WP���`"O:h�L�8��(ٷ ĸd���:�"O*ljčЇN�j��P���"�y�"ON�Ӈ1�(�6@�s��K�"O���a��L(�Ѳ-G(�N�7"O��J1
��%
��ᇌ�]�6-ҳ"O�軔�T6mD^����V).�� ��"OF��G��>�8<��ߢ
l�9G"O�A+�+�L`{�c����"O.��nX�b|̵A �J�N� ��"O1�!
�8R��E:A��\贔�q"O�K��C�8�\	���H�K8�j�"O�!Pu� Z4@*#�R��"O���Af��8PF�94�TU�E)�"O ���G !���qd�3�.�8�"O��"G�S�"����-��lk3"O�}j焍*.B$��ԯ�$��hɷ"O��H�[�;� C�O�7��ia "O8U% �.B��8�/Ս,��]A�"OR)����<pȾܡ�퉙r�h%�g"Op]sVH��e"���K�)u�$��"OF}��ޒ��4J4+�wc�T��"O�@�c�͸WԀ��d�6�AP"O��h���;��S�\/p����"O��K�<.��W�H�V�@i��"O��Ң�\NHֈɵL}q�6"O��U嚏P7���T�V�I܈�"O� �A(g�,k�=�@Ŗ$� �#�"O�ۧb���@�i�D�)��ո�"OF�Pc׬)�x8��F�� h"O� �5%M�o���]�88�"O̕�䑴fm>��b�T��&"O8L�E�?]J��P,v:e�B"O�`�R��|Ms �� ��<��"O� ��i�c@�*�NB�/� "�"O|ec���&ʱea�I
�1�y"NˁCQ����
�B ���J��yb�°)�%���k�ƕ��EF �y"�ޮ�zB���`��� �F˰=�K>!V�v�r���#O�8��Po��m!��C�Nu���I�2��T��둪X!򄆥u:�5cb-��x�B=+f�?K�!�V�U���ڷ�f�"�H�#B��!��"8�YB�k��
�&e��5e�!��Pܬq5��,?�D ��4T!���\i�bn��}��ݐ7aG�T<!�ڞڮ�P5b@�y�<y3A ��Q)!�d��n�̅��*_��� ���/4!�H�x����c�+F��ڧ��Y!�Q�B!*�J�H�	H�qEn]\R!�$�<�X�S��!&��)�p�۬V4!�.��`���Ѳ-��-@A۪^)��Z��H�����&�lr��V&�YLE�"O��(@���bJ ��P	 �>�1�IX�P�p���;����a��DS�AN"<Oj#<1��#&�f�Ã�ɿc�8, ��<y�́&�.�B���'�6�+q�z�<�c�A1>�* ��Q�c7P$j0�v<)��w�Mbn^�h�T�����8z�-�ȓK�zAxW`�� �����3��Ն�*_�ū���%��|jT���W��<���qNA�8>:�JW���^)V]��KQSj�W�
#@�k��=�ȓj�]�5��/;<8��n�<����Z�D ��iT�%��t�^/ZJ��ȓ[��u�F�P�$i���"e��^%���X�!���z��s����IL~�_f�Q� ю��ȱ���y2g�$t�|����l��m�a�N8�y��\�l?�H�@؍j�pC4�W�y"LS&疘Ц�;h����'ò��<A�'��'����;�zM�M�2���9�'�P��!�$��E␴!!�C�'%T����>lK�ժ$Z�	�'��	z�G�:v��p���	�ę��'�1�AD9j�2�הVZ9���)��<IB��37���a4�^}�<TQ��`�<�vl��N6��Q�)��)!��C�<��C�``1q�I����#	}�<9��>=���x���#z�<���H2g��yq1DB�(��L��v�'�ў�D�h���e�qB�*d �	�v<K$����b?�'��;�E	��}�� �&�4QO>ɏ��)�Ou���--^�u�Ã��^�!���k`\�VɎ:.�$Diޔ,�Ҡ.���O@\:c�Т�hG�p����gA8,�!��j�p8�Ώ�pZ����
'y��IM8����$��.6�52�b�!���s�-D���i͹:�<�&K�D$��p�,ғ�p<� ω�m��+���n��ap��V�<i���"���,��R���3z�<� ���5A�P�	Ё�	1�DI�#"O�c7���i����Фj��8@E"O��"�e�R K���f�(I b"O�;d�$v��"���}��"O�i�`�M5N�%��0�<H�"OĬ){(8�O�:(�г"Ov�Y��ͨB�c��	�(�R�kGBH<��^���!攣"h(xS�ńB�<1w��y����f�m{��K�b�|�<��G	�K� ��Eș2k�-��Xy�<ap"�TD���6J.�yㆯ�q�<����
!~�Eq���,9�T�PS-Gj�<Qf�|09����3t�������@�<%F��,�$L��ū��EX!bX�<yfbI�^h0T���cņ�k$��]�<�OF�qJ�CD�&3�[g�E�<� l)l��/6-����Up�C䉼]��41u�4���N�B�	"3FŠ@�ݾn_�(:O÷gD.C�ɧB���;���c�h�O@�H^JB䉧��l�FPp�|m�䠘�"�JC䉤I;��G�S�_d%���@�SK�C�!G'�鉖"�7Z���d��C䉛bA~�`P���V�"�P��̪
f�C䉭(@j���E�#� D,0�B�ii2�e�0��ՒR���F.���p"O�؉Rƛ�=��T,��i(ޤS6"OV�$�Ƿb����aZ6E�a�"O��p0ByZv��@d\0	��"O��U�J�7/ƝD��1ڦT�F"O�I',�O�abdP������"Oꈩ%O�G,*#�RW�H �T"O���f-E�G�&�`�G���A'"O"u��f��y#H58��\yRX��"O%x�)�������G�5qh��; "O���t@ >Oq�|q� �d�xQ�"O�S��A4h\+�U3:�� 	�"O�@�7���Xj�v>νzB"O$ܱu�E�`��p��Ä'��Pa"O=��p�0�r4鍶1���k"O���A�O,�X�Ȁ1L�R��'"O��(%,���.��a��{}:���"O��[���9Z�֙P'�,cL	Q "O�I�����l3p�U�1+p�"O������*Wo����&Ҫ(ҵ�t"O���"iJ�0Hp�G��C֐Qi�"O�L��B�������e͌Exf"OXeH�߀ylL�fo��g���"OV�pflD�j�� �-@�K��	��"O"�b�a<0X��#��]bV��P"O��Ǚ�$�1W*N�$-�q��"O !�2�Ĥ���C�铏>l�T"OtP��Y��\�q�t�Y	c"O����oڸ<=@��H��WZ��q"Oq�H�l@��q'�p3N}b�"O�Qq�>1P��c�,OJ+�"O2IIH�sn���E�3c^��U"OHAX�c�g�h;C�=nb"O�1 �i�]����(J+0�Q�"O����W�Cs\�U�-J��X�p"O�}���ՏQt�XZ��_C:��"O*t�Pa�/d:�!�l0*k�"O��ԍ�X�.�:!KI)�b��"O�Ī�H���UP��Y~ⴋ�"O� tP#��
&������B�_q�l��"O�e�A���%r���sih����"O���"D&'�$�A��=���Æ"O��@�!�K�r)У�4|� -I5"OD5��NM? ���tL�R�B1"O|�4�W�T�@h�Y<w��5�"O�p��qzD�
BK�l�t|�"O���S��)�r���J� ���b'"O��h^{9r,1�˘-��eQu"Ol(b���I�b�[��X8Z���0f"Oh���bG0kÚ嚵瀮`�~�Yr"O�L��f ��Y����T�V�"OpY;�E� �$�J@�ԃ'��q�"O���ɘ�J�.aҵ Q
_�k0"O(D⇘#k��q�]� C@U"V"O�Ĳ��-x�q�/đ[�Đ��"Op\�r�D�c
]��#�"e�~��"O�}ag���\: JB�ӊ&F8=�"O��#o9}1ؓ�G�)AJ]�"Oekwn��^�h�9�%GRt��"O���6a��'�� ��H$t<���"O��rrcő7t"g]1�T��"OFA���'��p�EA5I�@�"O�����? ^a��P�P38��"Ov�!�G�?/���E�V(�@�"O�R�?F�˃��(����&"O�l��e�{ر�b��$��4"OH��ѯ�=�����鉻A�m@�"OD�'��$/���i�
��?t�P�"O�� u�Z��<m���8jj�,��"O��D+́.hTaf!^�'c����"OҬ��_�Д��ꁳl\��	�"O~���V�T��hgɟ\�q�4"Op`��eǼs�,|�ǌ�$1�|!W�'�^�ISÈ0P�)�qa˔P+8{P⎢Fb�������e��X�6M/G�>	����c��}�ȓG��i�2�[a|� �V�C�U��-��e��HH2|�N�: �̦Y���ȓ(ElI�ʷx��pd���I�܄�u���&☇
X���!�W%��Q��4I��!h����69��1��Hφi��#h��PI���Ƙ4��l2�P9�ř�C��0��0x�� �ȓ#s��X��Q4��-�C�֧>��@�ȓu�i8瀐j���Å��GZ�a�ȓuǖ @RIL:1�ؐ;2mG.5�b͆ȓ;ras�j�?����M��&���P�0���ȇ�x���1onj݄�6~��@�';ܪ�-~�vd��x?q��.=R����:4�ن�/ n48e"����84fڄ{5���ȓ,�(�ٗ��9��!d�T� ���F����%�̩
�I@�_��x���M�(q:�+Š'v�Tqփ5���XyqD��t��`0��-� �ȓ5�PM;��3R��yh6��7��@�ȓ`&��%M�F��s �^@���P���F[�ra����ɝ3[B=��;8��E$0���U�j\��g:�E��(L\@ r�:_���ȓ)��gB�>L� ����4`z���dt̄�����E�%��W�(��{p$X��$]�ת�Y ��|Й��;����E޻o�p�`�	�b2�M��S�? 2�p��r^4��B�Q�p�Tqas"O�`[C�G#:F��QkY1�֙`B"O�5�9A�h�+��FE�X�8�"O�1h����bg��̕
P� ��"OD�z�i�=n`M�%�G4�n���"O65��ВH��Y����v��@�"O��b�nT�++��ҐMz��00D��h�g�",,�&�[;W��Ȩ��.D�H�uş�I����F"�(4�`e�!D�`�2$O�L�����z����2.9D� 1�*�P����P�J���"��:D���q$5H��=���[9�h}��=D�X�`�
�qBT+��#8\5�5g:D���b
b�9�5�|� hE�9D��P6kʽ>�p�b��G幷6D����B�!"RHx�D�JJ�H���6D��%��D���2���1���x�(4D��6Ɣ57|i���L��!��2D��C��P�_q�myP� >!ڢ��3D��s��B1%(�lB�d�#XKN@td<D�h��#E6$ �`���ܼp�2����;D�|���Z_gj1��� ��9D���P�B�a�&�T�Z�5[Ȝp�h+D��9S�	M��a�Ai��pQD)+DJ-D����a�#��]�Ơ=.s���.D�P+0�ۜ(d2�!ᤎ*
�m��-D���r���B/4���a�q����	)�
�#���s�#o�9��T�D&N��i:Cl,D�����.n��Z��O&�&5�%k�v`��5^�v����B0RS�&^{�9{@��f�:���I/=̚1+`MP2g�f�0���~�ԋbב�~E��r<��B�}y��"u������yR� 0����5ʍQ	�X�� �:��Q�T�����f`J"�����'u�Ό
4fQ6��MJ-CI�����,T�iS��$U�6lI�Od���I6�2�ʁ���D�E���R'�\Q��ӯ���i�`�O	5"�6�4���-�O�U�DnQ!�@�ݣ/���4oK*kS�r���zB�	�D����K�!Gπ|��¶�����<��4$�I�]�*t�W � ,����Sk�#Cǐ`�E
�~ ����L<<.:����M�l�����t���M���Z7//+�9bE&r`�aK�Cz��2 .�'�Vܳ��]�V?ɘg�\-�`*1�E<H��iS�#э{���>�vKL�p����F%8l���"�/o��ʰq� !1�`��[�z��e�8ޮ#�MВV����헚^��|�7	M:J E�MӋR!4�Q/������#�0���	����s�ۉ\`؊2k�/928`ə�4M���5���*�x�B����Y��ZXr�Ң���/7�� ��;��!�Ub8(x��`ϸ]�L,��VԘ�hr�֨N��q���u�ihE�K�&�r��hn�*27�P)����i�)�bm�F����JDJ�:��>�>tq�Ǌ)rڎ�"F�T8�,�e/��YK�J�Z� Z��زo6���DVJǦ�AI�-6\��VC�?H5fm��,�r��2s�k>���4��N�1Oh���j>P%�x;�!��p���)ה>�F��V	��!9��8��_�A���0 �T���;�C�Q�$#� C��Rh�7 �X�����04.�x�k��|��ӓs��!���H�B�`�C�-��\���Q�l�d��"�(8�r�ʵt��yaEMO�T��
B�*��d�pg_a�&n��<L�!��!Y�Y�xE��0��0�����Ȇ�H�M��zp�x#!V
�~ت�L؊'����'�6b	�pI�����bMA8yv�\s��W�j<Q`c`*���	��*��\Zwg),O�X"����r_��$��$�]:d��V�ތ�gI�)8� 1@��@!U@5k�;���ҳ��	 �h�B�Q�Ġ��I�k?A�OX�B����
ĩB�&�� �xBeЄ0J��Y��	]���C�=Y}X�_�l��5l��V򵃰�@�h��;K�(51ug���D�a�g3콻��Sv�����'*e�`(^]�J|s�Y�'��U2��4��5�4M��2럧 E��H_[�\TY�$،#��iR�B��
2~u�fEW..�ƉH�ヂ��Yr$��Ov��'���קjR�D��q�J�� H#��4�3n�nD,��N���+J"?�x�&��1u�\5�T��������JkupE1���-��}���K?Y��R��'�Dʗ�*�|}"4
L)XW����F])�jkR������«)l܉���2 F�����:(����2��
�~5+"� ��ĭ����%ܭn�����4��5�&n+}�M�Nn*I3`�]�s}�����B,]נؓ4�4��E	�Gʻ!��X�l
0|�B
�EɬEp��pb���7ż0�7)� Z��Z�'#�9����ߦ���\�xـb�d�UIp���2/��`�%�0qV���Ӱ�ZS��/[�x�`b�c0yj��GGz<����N�S�t���'�:�q���Z�p�OL�Y��*��E;F:,!I!��5����E�ީEUD�T�rӎ��1f^�;���k�K
u�z@r
� ��rѦ�N�h ��W��ʌ�e�'!<����[�BJ�B׳m�V��%��% =栛�˨bD��i/Y�vhj�n��a!�`M��$��Z�Ip�iw��V�|B�1S兾_J��'��$զO��2�e��e�5��8a����K�@\��	�aۥY����GZ�l*��KE%�60G�0�KUUp�ً&"H�PS}#CD�H�����H*�����!C�����^�|�*
��x"$aϬ�&���a�)���3�(W�@����ҟ�5�,R�,��"�g��@P�j/אxA�4MJ�c�6s<@Q���9X-����%4^\;��oPѺ�%у>Ypc�4t0Tq��U,9Y)���S<)�\�#6�
�48�FN�N
���ϓ�$���M���Vϊ��2,�[P|r��*j�1Y�ʐ[�88�3E�wIҤ.]ϐ<�@Ȭk�ϓ;��'GfaF'�Nu(4aC(	��=�J>icH��)�"�dw�d�L|rT�,#�rP�O�cs���`��/x�t�Eǵm��t)ښ�p>Q2���ty��(:+�x0gˈ�$����/W�~��+�∇s��D�'�v}�ߴ�?�`^��8�!ޜVΈi���Y��QsGG7D���7�B�uY\E�A��@�*ذ��h�$Q8�NK+	B2D�	�W��֟`�6�|2��.R'��A'�%l��̓6���0>I�F�4I&���0a�ZpR�o��9�e�A�W8�(O��/q1O�d��mF{	5@��p�6U��M>O��C���3$[��1�cW�����H* _!��`�D
��R��Q�QRWQ�<1`"��[8��[�#�i�J�ӷ��P�<�r�;3ŸB�	c�,O�PܓB��7�'�@*�
!Uy29��E�#�R%��'Y��pG�ӄp@t)
w���$$�LZ�E�Jܓ^$)Ê�D�\��S҇|�L�hQ�� ]��{��J≈ݚ0���\�K7L�3K��C�FЪ�9�=AWȁI\�vM�C�	����" �	Dّ�C,C�	�0�`���kC�4�6n��Lr��O�0������S����QE?��!�ІM�^T!�H?a���	v�=�z��JYD�,3�'n�R�c׽���`fڑV���	�'*���f 2��9�fV�=��}���Kh��ޓ5D���L�,T�s@݇PU!�������ƙ:��Z4/:W!��sʤS���������iS�0�!�č
<I�����`����i_5!�!�(MR^�C���)�.���eX|�!�d�5�衐f_>da�u���!�>
�2dXQ L�*�8(!��R@!��y�x����M.���4ϒ��!�D,��1h&��[�NI(Ќ��g�!�DJ�J����b̅�J�H�C�$�C�!�D�;M�\�T㒷��,IB�@�!�$B+:8�r ��&}�:�ևT�2�!��V�щ���o}�$B����!�$���+gDۭ&9T��u�J�!�d�%BK��J�!��P�<����O)!�D�4o�8`4E�>�¢E��!�$^p�  �"�)2kxAp��� Ρ�$��R�V�����!���;���/�ybI��R�Fqc�N�'{�	R��y�.�_lt=�bÈ�V��p(�$�y"�J�����k]�{�޽��M��yR�Y�I�jt
���8`��!�4�yb�� f"8��wě�O�l\��#S��yB�=b	@{���L���ٍ�y�"� p0�ڤ���)���Zۏ�yR��)n0h��덣,���BR���y���)0��4R�L��v0 x)!�� �yRk�1=�(�GE�d���`���y��{ri�)��T; �b�OJ1�y�'�iv�C0&ۣL���7����y��cJ%"=9��Q�C���y������0ì �j(x�kcF�"�y
� �!Ɇ�	BQ��I��	�%[f�I�"O��H�ANȽ+��U*,�F�	�"Of�����l�
t�M�i!
P*7"O���e���-��a�G�±U}J�$"O�� b߮d�x�dL�.<4J4"O(���V#~%�&a�a�����"O�[`*�;<�����!���ԙ��"O�Y`5��;2ʢ�p� ҡb(�f"O��բ !Sy�8ЯU�Zz9ɤ"O\P ��@��R$۳N�.e�"O����'{T"��Q�^�: "O�X�a�S�n�䑣�
�.s�*U"OZ$qK�3fH6#� �|b��w"O���+9-́���IQ ٨`"O"�{%��&X�y��J
Y�)@�"OL	���!�8�P'�$����"OZ��g�	
5J �R��w�p�x"Oni���Ƀ_�i1 ER�6�
9��"O����#f��J�%�b�8��"O�D���Q�gܚhR�Ċ1-�8�"Of�xd��H����%��'|�P��"O�<��D�)���sd�I˲�#"O�(���?*�ژ�)L&?��8B�"OUra��8I:�jt�K�^{�,��"OŃ7��-9��@�t�5��肱"Op,9d�ühI���%T�.�m�%"O�xx�퇺+�*�{��ƌ"�|X8e"O�.J�C��tJ3�3f2�c"Or�+!�\�S$\��¦��9""O�죀�M|��'��9 ���F"O䘉p��$# ��힖SK��3"O,;�'#<U�p	5�*4'۳�"O$����U��0S�#|�$k�"O�0G@X%Y���[�@�UgX���"O@YHUΈ�Q���3GO� m�q1$"O�6b�3~�q�V��F�UYR"O�yӧ�H$>�̑�MܰBr�Ё"O.A��B�9�U[��5(X�"OPU@� 1,.9�aJM�H��,�!���Q8�@S!W�j?"�4nH%4$!��8Q~݊T�B@�͙('!�$��N�ҒS�.�m:r�L�x!�V�VY@�#�9/o��Q�D��;!���g��MhG@%Px���b�@�!�dR#��E�H��W�#w�Şu�!�$������m��1��d��!�� �ܙr@$טj�~�#Q`��!�K�<p=�d,9�������#x!�
&���2KDh8@�F�� 6t!��]"R�%����k7����4j!�d����%b�p��phѣ�aT!�DS)�����C �#�j!�
2v=Մ_9C�,y�@�H�!���0+��;XU(�H�0�!� �qv��6� '}@YX�GO&'�!�d���5�Q("��h��Ӗ:�!�d�e�$�E�B	f-��cN�/�!��ΥE����K������4i#P�ȓ2tVp)�f�$�����4;:$�ȓN��݁#�ǳL�0��3
�̅ȓ7�Z�Т+2a.������7�p�ȓ;vޥrW�҃^r �B4�Pk���ȓmU@�����2TV��4J\����Ț����N�Yn�R�! #8���S�? �I �[n���G@�"[\`��"Of�ZR�s�`%��%'7��2�"O���Q��r��1��&_�8<��"Obx�qᛖ5�L���F	�6o��P"O(x�#�
��t��׆Z�E�V�
�"OP��%��k��c��O�t8�"O�u+�C_/=�赂��\�Q��j�"O0��&&^�����P��R"O�ͩ��!6n����7�ȹ��"O~��%�ـ(.�����P���� "O
L��c�"H� �����B�c"OZ�svM
�q�>�Ӣ/O&!�6t��"O=�r*DL
Z	Y&�ֹ9��\�&"O)��FN�;qv@���@�D	��p�"O�Bc��3�:�X�g]�@R�L��"O8Y(7�w|<,�f�8&�9�5"OZ�a7�.J!�ig�m�`��"O��{ "�Kΰ	A�G�}!�"O�-#�.w	�	cEH6�FT�2"O�e��?Z@`�C�N4�芓"O~�����hSl�s��O��Ȼ�"O��9f�ԯe����b��Q� ��"OvY��L�q?�*�I�C��"O� ��!��	r>h[�%'zHy�"O h���&Y��8�E�:���3"Olx�E'IФY'�O^�lp"O��5�=���ɍ�<fɓ�"O$@뤀)j���	ƦW,V� �Z�"O�}a�`�)�*XJ��P=�1�"O>�	���kX����Թ�"O��i��P�6&rd��"|�10A"O�m��
&Z-�Sb�}1x�ӗ"O�\��A9fH����G�;;:�a "O�����O2�i,�H$Du3f"O�囗` 3L�jPlF�b�W\m�<�Z!K�L̓0-��v�\��q��k�<Yv̙�cA(-Q������b�<�����l�.M�E��	>d��q�k�<�')�/%Wvi�cl�T���Z��L\�<1���r�0���V}�ȡlB�<�al_-KW%�U���&����J�F�<�r�Wv�a�*��^��b��<1�˕g�|��P�ࡒa�P�<!��m����EInN~��3	�L�<�f�]ZP:�2%���[U�:��O�<	��T�0p�Qc�Wk�V�6l�I�<�1�@�j�%�ŏ�YX���g~�<��/b����Ǌ]Y691��t�<!3k�5B�zy%�N b���WiIw�<Q��@�@ٲ�D�SL,�QLz�<�fO��Iu�� ��O%:= wB�l�<1���?\��L�v���Sʘ�b�i�<�r /P���NF�9LRr�B�e�<Y4d@�J~�ĩ쓣W����MO�<��a��1��S�;�*A�dc�q�<�W`
OtnT�0˘�3e<I	�lW�<9#j��^Ax����A9}0��R��KS�<q$�a�^�2u��7!��)@7�K�<�TbS'F�a0̝0|7�	Ф\x�<�S�P�B��E�3ʈ��0�7�Fv�<��eߵ���H��ܯx�.-1��^w�<ѴOs���\%��U� #�	�!�����L�0y�4�	��ɤ>�!��_�@����T�rt��HA���d�!�� �u(��0EX���CÊF&��"O�EѤ�,&ra����#�x�@"O2E`��H3�N���Z&z.l�"O���7�D�bR��P��I20�B"O�����$Kڕ
E�_���[�"O(��P;?����cFP��Q"O,���,L1(���B��o��5�E"Of�
R��QD<)$ V�(��"Ol,����2�"����^H8А"O~��"��20Dة��N'js�"O:а.E�P�;s��ixnu�""Oͨ��%�@5(t��A�r�"O�=[�G�h��@��$����JS"O�hj�h u���`��.s��L�d"O&p�2%��Z�Y(#'��s`$D�"O������ #@�0c�؜1t "O� ѱaU,3r����;S�X�D"O\��/��Ofn	+�m��H�:	"O��sP��c����� "�� X"O��"q��Wk|� ��C X`J���"O�EŎ��DƬ�C�K�Z.���"O"]B5�F/�h��TP�E"O$�@���)\���X��.�d!6"O���%PaP�5$D��:&�� "OX�I�-�I)���C��n�#"O�=B5È�)�cX+��"O>6�C�3��gA��d���"OJ]Iע�-](�uj  ��)Z��4"O�������C|��q��0O2V���"O<Q�BP�:,�0C:��X�"O�-�ŬK/��Q{SB�"�Mp"O4<IG#�7j����O�l��9��"Oȼ@cirr��㮕�P�K6"Ot���(+�`5���B34T(!"O��em�-\������z$���"O1JB�b<i�@ "m��S�"O�m�3aD�J� ��0,O!�@Xz��t��M�4�Q�L�E�!�DB.\U�Ȼ�Mژ��CC�_��!���B�tI���
u����C� W!�D�q�������Q��d��!8\!򄕧J�>X�F$h�pS�ͣN[!�^9_D�%0��J���G@�=m!�DȋW�P�qD��(M��b�&�gS!�dM<� �� �80���֏dH!�$��	�BB���>��x9#���<l!�$��H���`#Hٕ7�j%�TB�z5!�$�1��A��`��B��`!��!�D��p�3 �);�H�e]�5U!�ѱRU�?S*���	c"!�Ǹϊ��P���g���r琿W!�D�>	�x�2�$J5��� �ֺo�!���#�$�]F� z�pv����xXtK�6XDȰ9c�ςG��|��x�bI�H-Q��}!Bn�Jྡ��8���a��׎[��@a���	9d����*���B3/�f�U̃c�Z��B�XQq�I3,
� ыYP���ȓg��И��Io&2$!���"Z�ȓ;,��4�[P	j�H
�8�܅ȓ�x���Oԯ�\TPgDZ8J���ȓ1�Ѐ�%!ͤ	�����ݹ/����BIP(�5kBt91P�(S�s&Єȓ�]i5�߈2L��,�sq�y��S�? @XJ�)�4Nj��f&�(5����"O^i;�/�.�L�I��ܶ��r�"O8L;r$
Hq\��c���F�=Ò"O��@S�	���`0 ��e�jXR"O���v☒t�pxH �ѹ\V\�D"O�lh�L(�
�"�h�z��"O�l;��+i̅2�ȅ�L�^U؆"O�(OVk@�1�8H��"O�m!�K�pdP����E�����"O���Y�1m2��S�G�:��|��"O<�Ȣj�1>����i�,�,(�w"O�%H�'��!�080��Im˶"O�Ể�Q$�M��\�D���"O����Os��-r,�|�<��"O>\� � �/=б2[�g�t ��"OTl�q��r�VH���4Oz�l�6"O�q���u��*�*!�4��d"O��K3
�8��5\  E��"O���,��{�εc�c޾k���'"O\%昌S�ND�ʳ5!�"O"-*�B��;���Z�	48~p9�"O���Q��2nFx��ď���+�"O��c���[��L����vUp�"O�8R�,ĴD��2a�D�W��1�"O�	��O�(�@�!3g1Dɰ�"O��j祐9��]R&�;>����"O��(�F�L�]�=)��� F"O6,;,��b��	�iEQ�:��A"O�(�fc�:G%�b-�`�n�"O���A�,'�b�0T!N9۞���"O@ؐ���G�F��R �3e���ے"OT��U�S�V�v8k��վf��@�5"O��"G�G+-j��
�	z<��"O �R��9w�`�)I��I�E"O%!�i�F�X�5�Pg
|U��"O*8!��Ŷ��z�&O[��6"O�Pe��>!��(ȁU;�0��"O`���O��R�(*�ĝ-,�E"O\aI3#�)M�@ISR��6���"O��ٕ�	T�L���H��Ce"Of���%�C�ؘ #���q����"O�=�ł�L4`#5�:x\���'�V�St�_�Pm6��@�\���Ů�3"��R���K(�p�ȓQ>��T�@� ���C؄DX(8�ȓ��0)�]�6V���#��(�m�ȓbY<"��͒R�꼚E�Pr3|ȇ�5u�M�"`����p�h�E#Z��ȓ$z�A3"D6`�N��$a �d�ȓ$����'䃏T��h���	]Y�]�=�W��.����)Ա60( �2#��7D�ii"3f����-207�h�X����*�Ũ8��ҧ��#a�Y�T��!�*�97��.3�<
V�$�D��9y�q��'���@4� �]W��1��)�:i�A\��B��I�<oJ-��i�H��I��6Лv�K;��Y�ٍ�V7��z�lpas�T1��)�Z�~�S���<�^���	G2ߒ ����%���3˵<A��O�����5���3VA{���Y�����>a8�2����S�O���X��\4�X�Ï�#��!y�O�䪁�ݟ�-�C>��܄m< <2��Ǯl�nH��4���.l�l��>aU�X�T�H���*%5"�(�<Y���0>�Db֌JB%Z �-^f���`Xw�<�LwT���RWZ�	U�p�<ᗪ�r=i�CH�NP����F�<)@�'<�Q�fP�NSZ�S�
�C�<A��ĝ[� iM�4Q%�����E؟��>d��P�c\�~\��6*���S�? vL�㧖X��i�Oϕm=��"O~@�e_�{%֘h&��Q�`�t"O�)���$E� �� �HE��"O���OJ�>��እ�غ ܴa�"O�H�΢j&\	5i�!7�ъW"O��M�;z��y4/;�X�C�"O\�j�B��n�V@g�L'"��Q"O���uII�u��X#�hHs��`�"O
(�q%�BFd�ËP�H!�P"OL�7 �(8n�� ed��"O�����Nټ�9��\ v 4q�"OH�D���k���(1��R�"O�Jc&^�W@�g,_�UO�s�"O"`3V�^61��E鑄c>R���"O��8@�q�ɐ��^&n��"O DV�{�"��A�N�؜��"O�0SnQ�`
Pc'�]^����%"O��0Q̖$@z��ǁ�;[�%��"Oh3E��S���FV�g�`�j�"OlI�H_c|1JP��Y���K�"O��� .\�2���a�ΩC� ��"O�aV��D�ֱS�F�?%�ui�"O"��tA�8o(h��D#O�H�c�"OT:�c�� i��	/{HA��"Oة���:�x"㌻l��{3"O�-a"n�0������C��a�"O^�f�ފE�q�,JC�p���"O��IV hq.��(�3�V�P�"Of�re�Xr!��<��"OZi�-��{;��p�o���|���"O|ĉU�ߡLX ��NY��0�"O��!X�^��Q���Ⱦ2}�4��"OD�'�:w����@��F�Jj?!�dس_a�{w�L -��a
%!�D� E�����B�_vj@Y'��!���B���xrkqdF�rR���n!��W��)H�fL`8 ��~!��S]L�i$+	/Zi���\,WQ!��Q���M�3(�V��#�.%/!�
^Y�\h��j�H���ϩ,!�DI�3�0,�!@����#�a.~!�"�� ���	]��!�p�H�!�-V>M�E�C)~��(�$�Fd�!���K������0@ҙ e
GJ!��A�W���j�%#]�,A�U*�!�G�E�T�"��{�Ic��ѝs!��	vz�8PwhA;^��KQee!�D���(-�"����d�2�Y�!�dD>&�>8��*Ǧ �|���aHs!�$^6��`��Y�9�·C7!���MHsc)�42="��*�!��Ԡqyl���+�J.�$�ƨ�C�!�DQ� ��%K��+Q+�� F��V�!�$�7�y��
��D����R	/�!�d]�WΤȪ�MǢq�r����49D!�J�>d���K�V�-$�O�!��<w��xL .�ڤug��M!��ʦ2�sE���[���0�!��\�'��ɫw��9)̬C���!��A�[��Tkr-@
n
�̩���Ag!�$Ӎ#�����J�Npj`�ډ7a!�$�>0,��.�C�⨪��S�sW!�A��h#�B�Y�,��e��[A!�D��5�0�`S�=�\�R��N!�� ���Ǆ�U� E썽5��q�"O�4{FiOc',����d'jA�"OF��f ��� ��C���:�"O���!��9|�"i��[�C���a"Ov<0�N�S�>�SH�!T���[`"OP<�3�X #�Vt�qf%=�N�r"O��t��//V�	�D0+qV-�B"O�1)"D�|@��qD�Jf&�#"OHL3S���u�6������.�� "Op�DLBEʸP�'Π3
�2""OBh �bP�H���� �RH@p3"Ol��.-�4�2�-Q�O?��i�"O0�[Q�
E2.�< �'"�D�<��I�Y¶T�1/[����$D�}�<�jD>���S�L��>`"���c�<��g�Cfn�1�p�N!���U�<ѷ�]�
]:`�W�F�f��+
I�<)���-78��p�+}�hZD�<1D��� ��l��H� g8jB�~�<��N�<lZ��]��*[�I�O�<Y҇Ʌ{�<� ��m���H�p�<�c�Ը3��Maj�I�2=��O�i��hO�O[��P��b(�� ��;�'kT�!G��)�r����ٱ	u��{�'��p2E�@�'��TbC��	�P1!�'���E쌓qx4�,��&Hb�'��xKT������!G�j��'�)�SD����m��A��lJ	�'����hŚ���P�E%8T�
�'�bU�Cو}%6�1E#��x�Z��'`@q[���R���C��r7|b�'P�a�i Jw�=�$޿q�di�'�|� BC
B�yq�S�ل(x
�'�J-#�OQ�}�0I�f��N�@
�'��!�S0
1�i ��Z�_�H}�	�')�X=a�|�31�P�[�*k
�'�z��ǄB?�������9]�

�'�:a��F�E��(рǚ aA�)	�'���������XH��,�
l��[�'f&<�%�]�K/��C��UX���'H����(�&y����M<SOp���'0� �4ݍ��!Z�M��[�К
�'E�$�bg�V���ԥ[ %��r
�'H�J4�ʍ~��@�a� FD�r	�'�B��6+Y(ۖP��N���i��'9FI�6.ܨN�,���e�y��c�'�p!*r��=+��li��*P"���'�Ҩy1�S�#�X�8��دs�R��	�'t�HsC���|�`��#��a	�'��ڦ����K�l�<ETҹR�'��$;��  a��˒-ܫ0��[�'�ܐ��g��4)v�)��v�@1��'�&,)�mǽ�8��$
�W�`!;�'��E�Y���F¸�S���y�F_E�a ��W�����dՌ�y��V�. HP&B ���;1o�$�y�˵a��XVN(k��1�'���yR�ڿ>���0����vg\�l縴��+���,�{;܅ꖠ��A�݄�{��$z%$��x��)B�iLY��̈́�o����� �=<�b4r��Y���Ԇȓ&�.�IC��S&8����Dm��7��!�+�J7��ѳJLd��m��y������oR��P��	HE:`��S�? ��v����x�d�$9"��"O��;F��Q�]���D�`�X���"Ob���8=Қ-@��
�g��"O�9c�ƞ�L�B咷��dT�x[�"O`A!�V�m蠋 K��S`��A#"Ol�+�KL��T3� $/� �zA"O�0)"�
�q�����O7�rL	"O��8�&��O��麲�o��T�"OF��6�I"v�<�n
!x�"l8�"O@5�Bk�T�N؛����\���"O���ǌ+���if�B=v��5#A"O�qIō�#E�ð�ɋZ��y"O�T��RR�����$���"O�q��_1�&��É�PH@,�u"O �c���Yh�9���!`�lAR7"OZ�)���"a�L���	B�"O41�ũY�9;b��
��Z��Ec�"O剰M��v��x�مM�1j�"O.�ʵ��f�}�����-���"ORYK��%g���� (	։[�"O�d����<F�Yч��W��{�"O6�@D�ڈjiAp��-C# BD"OhTb2-��d��E��+܇F�3�"O\�[��89L���I p*q�f"OҰ!�M��M����8*���hf"Or9S���:�����`�2r�R��t"Ot����R)�2�SA�;2rɘ�"Oxy��9f�ei����G*�J�"OΡ����9��K�Ƌy��8"O�MI��(K��=�p.��l��s"O�Y�� ��>K@i��l.�lغ�"O�q����Lg<��+*mX�@:A"O��Z���q�(�r1��>P&p�"O �Wc�=y׶�cA�z�J�%"OĤ
a.���v}�%F�?;��,�F"Oֵ�g��5S���Sd�$X7���"O&8����,*��h�#H0|+�ɐ�"Oތ"f*�P����V��=q0,%ʰ"O漠ԃL�%]̅cs`�7@�"Oj��5l,���{�n޵n��(��"O�U���U/G鮔#(U�q��S"On�b��]"�$��	ΤlS���e"O�l��]�x�y��G�sb��"O-A1�T�m�J�(�1_�٘�"O�5 �,P�/+hH�M�3AS����"O��ر�_�KS���n�O��4�"O9����8kIRH���$3�F:�"O�t���R�'߮T��zG"O\Y���ʄF:$Q�r/ 	wq���"O��i��c��,趭Փ�x`G"O���Ǆ�&-�	�!�,R�Y��"O��fIݱ*�A"�
����"O�(� �X�|�P�p���+�65��"O8�����2 m�:vK��Pi����"O,�#��(�
E�K�m,�0�p"O, A�F��%�
T��8"O�ĸR�O�v�Z�H�����"O`T� I���	H�l��
�b=is"O��P�oL��0P2��Q�R x�"O*�:�,�@6֑r�
/�N�"Oh\1BI(^���^�Ӗ8x"ON��Ú�2r3C/ ��x�r"O`�c6�'ਰ6c����C"O� [	^_"��P ѷQ{,Y��"O� ⵡĊ��:ؾ�����F��x��"O@$�)3ՄA���.h-�芗"On�c�FM�I����x��sT"O�H#w��A�H�C�-I3
�I�"O`5;���9y�yj�:YJ� "O�Y�5#�3�bp�$�\;Z�^�pu"O��@$$��z��}RE��"Bꉱ#�'&BoD�m�Z b�'΂h�6y��g�2
��DB�������ǝ{�T�����ӧ��	�(=o����a_*TSr�#,�a}������hP���m��G��{����R����S�(�k>�"˓?B<�	�%���C-L|a�	��d���\��䓑?������	��%ڢ�Xr���9(V�H�ї9?џ�0��Ɋ�6�!�TQnI�s�Ma�$_�]�`��<���!|������'%JN!�p�ŽC���Wf�6g��S����{w��yB�'�ndJS���V�À�Ǎ2̲��b��|�4�'3�HO>q�eK v�,�)n��bc�q
�Z?ـ�`��X�4X
���6r���j��!�e���럄&?UlZ j1<m�ǀ��]�V��f��*LK�p������Ҏ=RF�X��I�I�T#d,���`Gz��|�#��O<6͝'���*w��0D-J8����|2���!\���I�O:��|�ڂ��~k�m���;��P@4��959ᧆ�;NB��\]��	͟�S�&��㟬�b�T�I�м����XY��ʗEc��0�fO�
-}腑2��"~n*���P'�����E����7�ނr@��'���$"|nڢW{2��Q6-ʙy��D��-����?QJ>y��dF�%X����	Y��� ��'1�牄Z���P���An>\��ȴ��;>�	E(� F����/O��׏�3	c���ҥB#df�D̓)'��"cʎ2�(؁�A���8�ɨ�(�Z
�-PL$!׭F�K�Ո"�J�z�y�A��O̠���\��(t
l����ʧ
j J6�;X�AIs`A���x�	"d�������d��Y?˓�?��OD����K�+9�g�=R�:Ǚ>Y�C��f�� Y�6�Ƒ4� �s�M.Jj��nMզ�$�h��-��4T� �čG/�NX	��Vy��3u��$�"�P��U�E�� ���F�<I��%��[����uGE�O�(��D4�d��3���°>i���v0�X'��Z�ߙ`��I� �K�}�B��QH��/��M���dCM��im���a�B� @�%е��%�\��ԆP��I�	ry��'��O�S:9�ݒWGA�Rj��v�x%F�;��D�A�O}Z��+L�Dc�a�s�N7M�iz�'�\ԩ�a{�����d�P8�?�K|�V�ӆ*��t�ۗ5羰�C��o->��D.��yb�'��ř��T;q��v9#tF��92��[�!ëy�RP�Eb���HO
	B D̔.���{æۥmGb�����|�C!@��mF��
61��a�'
iR��?��i2bV?i�կ��@E�!�_�]���>|4}�IA�S��?	F�¤2,��1E�˺0�|���Fy�+�S�t�?`�b�i��(H��[t�h8��F"z�T�ZM��m��<�N>�}�U� <  �