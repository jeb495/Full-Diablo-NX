MPQ    W�    h�  h                                                                                 !"O=�"�`�%���)�Ŝh0�A$�Lt��~�I�6�f�@YYA�Vu��!N?�7\<湼	1>c�Ko�-����Lg��J�lV�;"mE�;��?�Y�B*z�t9I�)��/���7�H%|��	��v�$�+p<h�qE�7k\ߧ��|��3�� ��e_&��?�NT��b�*�;��`w�i���F5�m�?z��xCc<&*��Dz?;=�%�ħ���K>�%B�s 5W���Z�X�{�P^�i��a�?�ZM�+����WnV\��s�&nF�}������L붞J�?�b\�!��.Η�isΪ��c��ue�X�m�Z���5�� C�ܵ�6J�XȐ,�D���_��".�NZl�-�gM"F��yJro���T$P��"�3:W8|�!�o�i�K��p�
3oX�?�0��2'U���N����E#��7��W��h��ۺ�73~�aM�D�؜(�'���Q��m�q������ZgZ�TV*�G~�#.b
r��;0�s;L=�
���O�lYd�h���Q�~^��@�Eu����K��)��t�����) �BE"n��1;j�M;�dG�,��A)�R�i�JpL�Y�����"����1"��@/P⾰�Vm���j<��͞窰o���J�>T.L�53�řg�[dkά�����&�w?5*�V�Q(ӭU�"/3�E��TB�^�ms�	����?�L��.�da�àc)�пr*������\_�$��j���8��c*��n�3@�=�����ܟ�	ς������)˸N����6�֜�E�@X�uW�85+n�����Ƚ;^���B��f\����W��{�~�|T�L�����\��1Ze��r��n��ç���ME)���6����h�t�jV�����������F����ɚ������o�>/Ü|�Ծ�d��V��ŉ˜Z�YY�4U�52��pJ�ǌ�W7�T�[�٪��h�t�@�cvBނ����!�i�U�b��P�ֶ�-�xɘ��ߺ�G�9�
��T�nެU��.��4aR}�}�J��
ʹ"�d1V]WE%�3�x�z|@d6��\�n����wiO7mx*����/1�P��,gz�o���tq,$�)�Nܛ��9�U�U%5�������M\�<Ǒw/��>yiZa�&y����)��⥫>
A=7IP�'U��ȃfn<7(�u���=|�����3BjZ\O����x�!-��P�C�K�T OҐdie�������2P?����(Ȓ�}ʥ
�}Fh�3��(]#㦛:�>��2 �	s���ɴ��Vܷ�Q4X�Ƕ�6�O�U����������X2�
 ��O*��h��
G�$���?��sv�M��U�f�0� ��~o@�z�@�MKC�ݧ��v�u1���iu_�D������ݒ�al�~j�wʂ.�Sĸ�G����|(�E#��7Kx���z���-����6�1��tOVK���Z~��r��#����e�N�(��k�#���fx0ԙlH/�yDz��B\ �Z�e\�n�b�)�kxa��L��x}n�Pї R�=�G�	�D�@���>./��ƹ�ሬ|��$3Wᢍ&�'dѭ����>���q#����(�GGz��L2�"t,�g�
C�A�[�bPg=(�D*u�����yZ��pނXh� ��`��ӡ�s/�B����<?���t���I��eHa�����3��
WB�L�8�?#`���jr��(Y�� #$�=T���JQx��`I�W�m�v�h 88&��&�`�v� �7���l����C�!�B�=���� �ʫ��ɺ�$��{����K��B�+� SI��W�n�$���)��H8* B�
�NLD�xG����@u�#���2��D5�PƗ?��w;���c�݈¢+P��D����C1�<�.�������T�������ueb|��+���n&��k��d[H̷peF�N�ĸQ�v�i����N���E1�|�b�z�gْǷ@�s\����ѣ�����ް^xB���ˊ�D�==��ђ���f��2�E�3�!C����^��S�F[U��;vW��-����}�T�F RCʒjRl&�Y�m�v��{g����N�pm�`&u b�ň �v�?+>����>.ǅ֚y����DYg��x6�}tܡ��79N��فf��K�,��*��B�d��G�_w_*S+fm�\4�`�ko8{6�:����
�����+�JWf�1�kp!�X�6??0c��*Lz��h� &7?�Y/�u�2���x{��9�\=IO��@+��Pz�
J8�
ع��������a�^�pB��m.���U|H�����7m�X�Iq[$ FS|�c����<1���M]������"���"�i4;r'��V�6&R�����<���*����9)h�Hv�ƙ�N^w�e ����8���p"���U��ӑT2��69U	�h�%7�������"����A\��I��ۦ��*I����J��f��u����b 0`���.6&�*����km���7Dz��ӧԃ�+,�(���$��	��mo��B������%�NkY��[�����=��A�������o}Mn ��Q�P��v	N��h�80<C:@���jvnZ�(�A^��q�V/�#V��d$�+bJ�+z;ּd7��,�v�h��k���ep�;Vr�Z�%�W�ZbF�y��NM1x更����Hw<w|�F����aܜE�^��%L�����<Q{�:�6R�C��X��q�cj̃�}b�p�]�H q�J�@F�3f��OG��R&�Sj�b �t�L���O�R8*y\�(�%f6��iD�������;*Ɂ�l�f�_�DW;f�6��p�H;� ���"���V:qN�q�����L��1D�Xv���BA'�`���]4�����z�B}yAk.~]�;����i����D���7�=�j�bsG	 y��Ajr�:^9��.:I�!wX$e@�H��n��0�dX��:��"r�5}��ϔdOi����5�-7��b��vQ��w�V�u�,:�}�������]7�rŜ��|
!b6Q0m]��$�F���<#{��_��Q���p�n <����1��p���Tx���.ӲYXs�IX�o/ÉR����D����k̪���]����A��W�3���s�K�kS�G���`~S�d�\6~�[�uz���H�%7Zt�$�rqeԊDm�̏���p�������ka��z�0+b��<!52�ѕ�����^�x���0��+��|�VlV��D�R�n�I-~nA���V�B�Ga�L�Ji�Ab7毤�X&�y}�s�O�¾Q�050X�4qZJ}}/�;BӸw� 6��γ����)�oM_���.��(lP���-F�Yy�k�q��$k[!"it�:2[�|3mDo��K�Ё�e��X��I0� �2��w���H���_��@@�Ҧ�sMh��u��V�7�T�<�nDVל�*��.�Q��m��%����p|�5d�T��&G�q�#)ɓr��0<��g�E
�o�*�DY��hQ-���o~�?�@��[��?�faL�d �t��x��)[�8Eݕ@�LZ8ҀO��?��,�l^��d�J��Y�J �3�c�ip]����1]{�@��ܾ��Vȃ���{����%Iu��v�y��L]@��������4���쪘��R�e����KӨ~�"�\k�g�`� �����m�p:	#�K [�G�H.�ם�~�cDx���ݎl*w̗#�$6�䦴���0f�hk�Nᯂ��5�m�&�ڀ}����kN�P� �		����Q�Ek?���O���V�n��;����x��;y�:��	�f7J���<
�.�~�����;�ͺ�R\�S�Z�zfr�0p�X��V�H0�B=��1oh���jѦ����s�d+�F�C%�$�z�����o��>
n*|�����wV�}�&=(�'4p��2jJ�Ԍ�h���p[�cy����he�p@�q�BYTH�h�'����5�K���S$cx�ZA���AGuVo�-?T!����.�ݫa���}v���_
H�"��xdl�W��83�C��g�@��+O�L����Li�t�x���a����P�e��G!^]m��!,,_:��+��T�9<�3U�"�䱇��)��(��<��/1��twxZ�nl���<�(G��AAx� PGM�ʡ�f�4Z(�y���>�L�Ʋ���\���z����-R?�^2y��))�k�����1��g2��=��xȭ�� n}!lnx(��_��t�>ac �.Is�D�Dt���Q��e�4�}���k�q�̄s�'ɒ�w�����E�8��f$�cg�
�\��|�o��������U�
��k�� �\~j��_ŋ��~K^��D��v�%��H�����?4"��=�M��l���jwc��	,t��Xs�S�����sU�V��x�Wzzx�>-o���q�a�q]wVF������-��#�j�L�N��팦�2�H�fs�ƙ��z����D�N�B�̅Zd�y���+���sks�座j�x8k@P�+�R0U"ǡ���:$Y.*W��,�g9�?�.W\�&���d�_�=V�>�ɱq~��i;�b��?��2�
�tgg=BC�y��٘P"�=(�/*����܎y��K�I�u�{2R`�-Ӽ�,/t����]�<z�L�fJ�B�I=��e��6���0�
2��L-R?��B�ۍj�X.(� >:!�-µ���Q��q`�c��	�v�f�8�A�j����]���l����>�!l�=�y���&[��$��MGB��F�!B�< )V�r�Uڇރ�j��)��b8���Q�Na�E�'��T�߻��Qb�m=6D�D8ƒ������O����5r���B���Оl�ׁ����|���uD��p�_25e=�����ۯ�	�4&��螟g[c�0��K;�)҉���M{@���ѩ��� ȼ|��:z.���,Ԯ�(�p���/�A&���#��6ъ?�q=�~�<XT�h�f(��f�z� �D3 f��#I�^\vc���[�Y�vR���asź��T�u�R��jj-� ��?��;�{b��x��+0`A�qb'#����z�_��K?>)j���:�j���Idgc��6��]tU�̪Q'N�2��o�Ɲ|$�,׼y*V;B��Մ�kw���S&�>����`E�r8�:�b�������L���E[�xp�z��Q�y?��ڊ/L����"7&2�Y^�uF�~�=9���[�y\x�&Ok��+�<#z��o8g��U������caI�p�sB�h��+Z�HVK��j�¹�$+�$[;F|d H����1U��M���aڝY���4vr�'$���1mRMs�����W���+ԝӕ.9ds�H���Ɣ��^�V� ��F�À��R�޾wO���T̈́��1��	T�%�f���M˲M��ʨ<�|}Q��5Vۡ*��{����Ą��ɾu��l² �>��8�6���a��k��(ǲp7�ҏ
Ծ5�,>G箽�I�Z;Z��ɘ���\�[6�䉭׭g󳅀W�,���I�9���&2�M���'�����v�88�����CU
O�x'n5���|�����Q�<�iաս��d?f-b��czl�����~���q
��ia��>:�p��\r>�q%�Ά���W��6NH��������*w�jZF�Č�B��7��^�X���`���g<l�>:�ʦR�u���܂�W}�ceK���Hp���H;�uJ^ũ�z��ߝ�E�>&�������/�~�<%O���$\�K����6��i�ш��(��F�]��*���l��_8��;aۀ�OP�H�5 �"���1q�b��~�����r��NX����O�'�p����r4�fM�Q�4=�AA�cU]��������4eGwenD��7!�!eRRbΧ� 4M@�\M������\DQI�pX�]t�C��ncC�0�[���՞�	�p�>lī}d�}m�����H5��Y�"�t�?��Q{VG���f�pH6:U_�������s���L����!�(�0E�����FB �E�O{�eיB���P��<�,쾬i��+�-��ٜo����렲4�����
�ÄU���������Ī-��]ʞ��2��Y
��)}���QSʗ`�1�j~.C���T�4A=�p_�j�����t�_�r���������Mۛ�<�zN��qɖ�KQ��u&n5������E�^��R������+���ѠV��;���=��S5n<|Y��^��L!��J��bU.��r��s������$�X �Z�G�XI��v�w��O6��i����A�_y�n.l�'l�q�ĝ��F<�y Ǧ�,�v$�5"��a:��|n�)o%�9K��n���2XmA0��Z2�-���$Q.�{~�����0h|������7)K���D��i�^�����QWQ�m^�<������cT�"XG>�1#$PYro]h0������
}�F��Yڧ�h����]~�R@^�&����8���]����t'p��� �)�C.E����g����q���,2�_iG�_�+J&͇��N(����G�h�1�3$@e����GV#�2H��2ش�G��>���L�jλuv6�X���@����-n�V���3�ӣǅ"��#�"&�#"�T�mӎU	^��� ��B��.:kz�9~Ac_NF�h=�G�����$�[�����ً�a�#���i���3���H[@�p�ϸ{H��O�����|� 0:����EF^
�+JM�n��n�Q�Y��3�3;��|�8�f���A���ک~��^�{�u��\�՚Z[@rk�����O���$�C;��z���n�h�.jL����������F�7��T�5c�0�on�>�8(|&�ԚV�����u���,4��2��J�{p���2�[��5�Q��h �@ҟ2B�E �C	ޑ�T����EF؎��:�x?<���!G�R���T\�R����.��~a�/}1#(�h
ã"�u�d�ڻW{83k��0Լ@���<d9��2i��kx9��&���?�PQ��b��؊ ��,�n~����Ϸ�9��U�0��L���l�,9<=X�/�h�o��Z\6�����77��ۗ�adhA�lP���Ś�f$M�(k� ��S	���*ƍ�m�L�\�B���>3.%p-�k�y�κJs/�F6X۪�%���2���e(��Ȏlʛx}��O��8(�4���?>k�s ��lsn�ϿS垀�t�-�4�o���̷����.n!���ت�,/�j�߅�0�^W@
�K0�7wàշl�C^}U�/��F� L$	~eY����ض��Ky���Tv{�Z��PC���:�X�s
E�|�l�rj�n<���./��N�������Tx�Jz�S�-J��ɬg%�f�VA�-��"����#�H�ǈ�N~�����䷻�fn���"����|TD��BR�uZ?=g��ȏ_��kn���\7x�P�wR����*t�����m�.%���o�w�"���Z9�Wׇ�&���dG�A��
�>�Lq�O��$n};w�V�2��-t�'Xg�$2C�m�LP�y�(,*k�ݷ��yаވ�ә�]���V`dv���K�/����0Q<�� �@Y���I�r-e����Q	�)�?
vLh��?Y��O1j(L@(�|� Yp}3'��zQ��`/���nvE��8��L�\�GWֶ1%+Ul2�1�9�!_��=`���.�ʡ�o���$6T��s�A��BG�� �(�؍����эE��)N�8`�� �,N�j n,��6��67m��&�쨭�Dk��ƍ�H�-�<
�ɤ�!����p���rdT���nܿ��E��("����e��BAI)I���&;2�Y��[~?��fR<����.T��3/��T���N�~%| _�z�ꏒ}����t4�������˰��Ȉ���]n=��w���9�f�w��%�����3ʇ��0x^7Mc���V���dvM�|��-��uT�ĬR9�jP���Ο���{]����̪���`\Ɋb��]ֽ汵���2N>$-��P+;�%A�n7g�i6r��tR(��E��N������7�,���*��B�Jb��I%wU��S!��p` S�8�:�N���)�����3-�@����$p��6�l��?&�l�c�L�������&-��Y���uF��Bq�6!�\���Os�+��QzY�u8"4�\��Wų�,aIS�p<��c���~�H���!f�vM���c$�PM|��1���1�&M�5�#��/��k�4���'���LpR��^LN��rq��K���Ű9���HM{�Ə�r^-�� �-X���2��'��R*Q�C  Th�>�,{�	��l%�B����olʃ�4��F���ۜ�^*���}9Y��ºʌu�%���V f���"6�Ѭ���k���-�@��k=���t,م@����ᵌ���F��5!T���a�6������H��]\^������T�e���M����b����v�}\��&Ю5sCp������na���.TR_�L��ħ-�x��dZ;�b@Rhz���ů�=�lH���^����tpћKr��8%�&��^�ЯAnNC#��Q���H;UE��wy�F{���}���Ҧ�^�,-��ҧ�jQ�<���:$CR���������c`��3?opC��HVS5J�iY��[�F�Ȩ�_�&�5�S��a��!��O}ϡ���\Kqc�[�6�+i��^�d�*��`� �*u�lр_��o;\�f��O'H�� �\3"��Nq�2C��������x}X�A��}C'�@��hi�4!BN���P8��A!��]f ��`ꯀ�R�DL�7�x�`��b)(z ��H�wP��0�7z�IJ��XZv��>�Xn��0FrH���+��e������d�����cP��5pQ@�=�/;��,,��&����k
�:�`�P"����h4i�j�d!�:�0�����?F�L] ��{�g��@�v�@��:�<&�[���S����������w��R���?��@�x�?��кd~��U�����]�ֵ�m�g��F���*}��&�S����'�~	&X�Ғ��F�k����bd���tߺ�rg�i��h��4㿦�������Q��,8��f���/�5�6��7��L!�^����r S���0+�4!�L�>V����G���Dn7�Q�fY��J}L<�J_�
b�㜤S�����s���t:��4NX#OZ@2�3�(��0���6��u�i�i�]?�3y_�Ֆ.G�Vl���8�lF�vy[�"���m$��"_U�:�Z|�cco��K�<8��$X(�J0ؐ�2�W��S��_�p��r�
X�h��h7����7�a��D�(�������<Q���mf��2��fy�e�T�=Gٸ�#�Zr��0��x�
�7i��?eY_h�Ju�G�~o��@|ճ(Z\0�ޤD�ڄ�t�y��]�) $ESE�Ԃ�l�v������,m����%�Z��J���D�ir��_kޕC��1��@ �����V~���ƋMl���_&e�L��Aζ�x�	�%3���|������2�D��"�Ӟ0Q"@M\�ݠo�>��ω�m�� 	���A'�=�.�����TczD����\�"����$l灦��8���ޞȄ������{�#�)�P��Sr��߫���R3��גG+QE!�K�fd��	�gn����H��^�;�EF��f����3g�L�_~�<α]�j�0I�\xKZ�%DrF:��.䧌?�>f��6
�)��h �lj��}���<@ȚPqF�%��Z��a��Go��3>�#�|aG��5��V�����C����4�Vs2�gJq��T��^�[�[��׾h�x#@���BOW��JD��Ġ3�?A/Ŷ	q�x�=��0JGk���T�Dˬ&1n.��acAC}쐢C��
>K�"�d�LYW�W3�WM��`�@��)��PͩV'i O	x�7��ݨ�@��P�W�}�S���}�1,����+�:�9�KUV^���1g�}�����<x�/gc�j��Zri`WC����v�ԥ<�?A�+P}������f� (&᪛���BU�h����\ 2��"����-ȼo��^L���a�!��_K�J����2a��� �e��P���}��[�q�(.�`��H>Ƴd H�ts/���:Sy�[È�h�*4)���	RJ�'�iBD��I��*ƪl���?�� @ջYgt
X[���q;��	䢾��Uzt���&� ��~`4�n�q�K��:5�vV�g��;�:��5`k��o��Ì1l.Hjm�ׂ�A�i%'������o��VtF�̪�x^�zn��-%!B��h}ا�V<��kP'��	�#G�BJ�NY���l�RO=fi�`�}�R�M.�D� (B�űZ�$��9���Ckiw��]m�x���P"��R&�?�q���6�p��. q:����s��u��WR*t&d}�d��7�s�l>�y�q4�����t���5D�2}$�t�_�gsd�C��l��P�W(G��*��>ݒ��y�ňA~i�"�1��`ߦ���W/jmH�v#;<�=)��U��oI�Z;eyܝ�lt>򤭖
軦L���?�����j�_�(��� t��@��U_Q)m4`���)v���8i�ūwYW��9֑%Tf�bl�I��4/!��=F�IE���@�Z7�$q��}�}�<x)B��= �Hxب���}��� ,�)O��8�E3���%N*�U�9�߱|k�����=MDT/ƈ��������.�)�����.`�F���g���k���؅֩�� �U�xe��f}�=�ڎ��&�X���[���xI�ߝ]�i�G6��@q�_fn�vU2|bz$\-�X:�$1�Ǧ^O��V2��2b��=2�*I��5�=�ioٲ�S�ԥ�fp���vv�36NƏ8�^DS��qE�
.vHi�>_�0�9T4OR�a�j���
��G$�{X�i�.䈈�/`w#Lb>J�
g���?��
>@֫m|��΃۳�gYR 6M�t�����N�n��%N���5F,��*LJ�Bv�^��G�w�OTSqբm�h`��8�'�:�]�w�6�r��]�;�^�B�qpR���g?�_X�\IL+���99&(Y��u��� ��|�L\�_O�y+���z��[8�xd)�-_eŎH�a�}�p�6[�^�K����H��/�<-��������$хh|�����x�1��M�z���ړ$���4��'Z9��/R�4@�������9���H�-_Ɗ��^��� N�͓�pV�H��-%w�~v�T���'L	
�z%h>ʹ3Z�CF&�^h)���'�ۗ-�*Z�O�8���� ���u�v98k_ �1����67���Jk�.yǨ)���g@�4�,t�������I㗌PUy���-�d���C��ڊ�{Z���m�r���o����M��静��!֗v�E�^��i�DC�����n�]1��������G������3$du0�b��8z̛�����쪋g���|٘���p�{"r4��%�T5���J��N>L��-���`x�w���FV�h��V�m�^� ��6F��%0o<�=::��R����3Eh���Ec[�����Up�:�Hq�<JT.U��Й�]Ǩ{�&��$�s�V��<4.O�����L\�Ko���6��oiU�4����S[�*ZlY�t_n��;W��o�HP�$ ���"|JP��.q�"����#�ݭ�B�.XO׀�!�p'x1��Ci�4\=���BE3?gA|.$]!!��N��*�}-�oD���7WFG[4'b��� �����s����H��/I�� X��$�99Dn�0�6�����6���:�kd ����l���5+��X�2�
X������H���f�]:� �o��/�"���E!�!m50>Ȯ��TF��(�c�{�6׏�
�Q�@�x�<��c��9X��v4=v���F���@���������@��z�|�3��uR�����#G]�.���!y�_��	�W����|�JS �s�'��~�(z��Hjl��f�H� [2�V�tt�5�r�F��U�@�q�ANz��9��0u��������kY�5Ï��F�u��^}e���n��F�+�߇�i�V����X��n2Х�g�4�x��LW�J�}�bȒ�����J��s�����ޝ�ad�X6J�Z�<M�ɩ���H�u6����ĕ���VF_o+k."��l����+�FRy��ޕ�5�$��"���:�
�|��o[��K�ݚvwX���0�xT2C]�`�ځ��'��Y };���wh�H��&p�7��ͤ,D�J�����¬Q(m�LV�(���,��TB��Gt�#��r%��0mz��!
sؽ���YP6Xh"	D��N~�Sd@�xh�C�L�G��K�g�t]��ź�)lE�Tԝw������N�,��,�r��U�!J��C�"M���+��!�=18@����YV���!ҋhb���N�:.�*�]L. Lα�I�YPNr�!��	�N��JgS�����ә�"����T=�YA"�J�m�*<	Ԟ����8qk.����c�Z\�^�ގ���H0�$�������A����hĄ��6�)Đ����܋����ܫ��d�a�:�ΐ6�ݒE��|ᡞ�{lnܛ�qsȩ>[;���.ْf�Ӥn���瓭~��ٱ�Y��볨\,:�ZQ+�r!	��'i�9�5�0�А�vhi�jB8�wI��w���5F�%��50���MA�o��>�.t|����к3V��$�7ޑ�E��4��B2��'JL�Y��\h�l[��Ih��@\�Bʈ����Z�U-����q<�7�d�fx�_��K_�G�k�v�T�����K.�C9a��6}�=^��
��"�Xd��W��3�d����@PUI�X�Z$�̈́�,i;�xo|����6���GP�M�Ø��%3�X�|,�����Q��9M��U���7������{ <���/~�ea�Z͖����������
�A)p_P~2λ�f���(�D������J��C��V��\����&��?-����$�@f����Q3r[���ؔ92�8Q������{ʑ�o}�78Q6(�}妇�>!�5 �`sJ�Qϵry�6Ҍܣİ4Ĳ���邠?��*�d\j���?�G�l��4v߻��T�D
���ȭ�נ|�9��UU�V�') �3~[/pt?�,��K�|r��5�v1�Ĵ�F��Ў0&Z�)�s�~��l!vj��^���uĤ;��$�k�� ��$���fmx �Tz�``- �A�"�i�B�V7k��+̰^P�#e
�+NN4���Wޗ���fd�ء޵ �D�	�BH�9Z����Z�~���/kdi!���3xi!1P=��R�[��؞�0q�ax..�%K��[Q���QW��&?��d�"B���>�Uq�>ʍ�3	���Q42X��t��g�:C�h��ǐ�PSU�(bY*a1B�mf]yFW��HĞ�j�`�g�l�/���Q6�<+�Ŕ7����INc�e4����o���
�ygL�]�?�"����jޒD(E�` �<�)z�0ȳQd�#`�&�����v�!�8$���90h�l9S�Dlh� �/y�!��=�͂�d��ʗi}�5�d$�h}���7��B�<� ?����:������ )�x*8��^����Nr	Gv㡃[��,���0���&D�?ƃ+��㤴�d@�I�1�R������p降����"$'d�@�r� �����e�gj���$d��_r&���ς�[�厷\�b����Ĥ��U��LoѺ�-�1L�|6�1z����3��_h�A�>��-�R鸰J�_�E����K=�՟���ot�f���wȔ�1��3Q�l��_^�Z3�2d(�*DovCuѩ�&���qT+�yR/�;j���E׀���p{S�ʉ��\8�`���b����w�+���h�>������|1�6g�Z�6(��t�.��{aN�<ȁ�ۤ��n7,(M
*ǝ�BQ�˄3f�w�5�S
���U�`v��8�b�:�k��v�o�q�c�i��6'?��g^p���?Ipku^Lfζ����&#;�Yo��uw��-,g�7�n\)R�O<��+���z0"8���D�g����i��a��}pr��Y��<')H��ǻW�l���$ۗ|5�����1f%MI��9�o�:����4'3d'�����R^B��9������r�d��9UMH� �ƅ�^� 	/��b��^��@���>T��V�"=�	e�%#Z�N����<��9.�-�����vے�G*�$*��f���?-�ug�'s� ����m6�~/����kٗ��#�7�c��o�,c���p��k����m�k��v�e��*P�:4��~Ċ�vw�o�-�e���_��9�Mru���F{��*�v�-xIF��$�:C�(g��`Cn�z��-�����B;	�z���^�d�E�b6��z�cļP�ʯO��b$��z��o�p|�r���%�Ǵ�F�D��L�N9����E��r{c�w��jF1����/��P^�4ۑ����.�<��:�6 RjpA�n)�(`�cV�F���p��H���J����u��L����&�;p����`kl�W��Os����\�Eo��W�6��Vi��
�ڧW�1���*5�El��|_	7�;R;�`��H&� Ar"�4���q:3�O�p�ظ��- X
���<7f'�A$���4�XL�"�.�A��]�a��.����f�D��7�3�VՋb߈� eP������&8���E�I�&�X���4�Knt��0��ȣ) ��z(uΡ@�u qd�h���+���5��Y�s�}����~G�����a�{:f�����@�J���^#� �!N�i0ٱ�����FS�v[�{ӎ�
Z`�,�P�Z��<\������<������ �m���˩�5�\�����u�����0`��^��i�][�����*:��+�:��78]SHٯ�n�~�K�Ho�G�a���{s���t�+r]�/���]�{&����훑��ꋸ)��uꀜ�s��]5��с?���8�^x���(�u�.�+ ��B��VZ� �>f�쵇kn-*V��x�3��LrC�JU]�b�aJ��A���s�#��*���|XQ�MZ6gy�V{�'Wݸ�Dm6���ː�Ե-xE_��.��Dl<Rg�n�F�y�ڕ]�($�!"U��:�ڝ|��o�&K�(_��M)X���0��2�N��;)���sR�L��x�Φu�h�Ģ�Ac�7�����6DB˙�/���8Qh�)m�SY�C�h�\B���T}�%G��#�r�PL0(`��
�𒽖�Y�-�h��j��Q~%E�@��߳^P�R��Zr}Pi�t����7�)�8E�tԸ��l��� �,��0'��P0J7C��U���fi�U�����1I@6���� �V4��y�!���2�넶V�e�{Lɪ.ά�}.���5����S�¾Q�	�X�Ӕb�"��M�S(��t������md�	����S�3�Y.K���j:gc��#��Ɍ��̃t�$�^����dٜ���TR�������vm����ω�*���y��X���N�Q�K�=*DE�z����d�?�n�p�j��d>�;�r����f�1��w����~�\����ͦ>�\G�Z�P�r��V�D﨧����4ҋ�א��Vh66jj��*R�T������lF�[�ސ%{�f�Y"�^o�@5>vY�|�3��k�V��2���_� �V4�|2���J'�������F[���bNshQ�f@#�yBE�0��+!���=�i�7=涿=�xp�i�f�rGa�QKTs8�\.�.�� ad
}b
Ny_�
4�	"Z��dX�pWL�W3��G�A�@���3�V"�_:Biv��x
�z��`��ŰP�0CóI~I�>�3�,Kg��U�K��:9��cU���\�s���S\<�q`/��C`�Z(�������l���>AdNP�#�ζE$f5V�(��K���8����g���\V���J�?��->�c��
���K��`��'M�!��Ӄ�2��b�����]}���ZPs(dd¦���>|�� �1seB&�0������*4_���;�����Ŕ[�E�"Z#�1J�V��O�
ڲ�hǗ�&ˢ�~�U0^K�WG� ;\~VJm��P��s�K��˧0VBv%r�4r@p��+%�����9l<ެjcQ҂u�V��q�����ӱ���7�BB�x;�zd�-���]����?V2��!'���#7�{8-�Nݱ��*w�֖f_S�3�*���zD3�B�>Z�p��6��0tk_{���x$�IPX��R�(�_�kt���
s.^ƀ�Y�Sc���mWH�&��d��`���>���q���U��Ι�+\23�&tS0xg�CSC�۲�"c�Ps�(}.R*ܩ�H�y�ڐ�w3�NA��g�`���(,#/`��,i_<f:֔���ߦMI���e�#������h
�W�L�<?*��k�j9�6( Y� �҂��V�QQ���`PR���GvV��8�V��;d����Gm"���lWl�*�p!pQb=�������Y&��+$�" ����2�!BX? ����@B�s��Z)�=�81�!���N��1��:�Aߧgl�je��Y�4D<��~�\�>��;��d*��"Ѻ��/��K��C����w|F�����ѲK�le����j�����)&L9���[����%����q���8}���x������b8|Q�)z��ܺԚ	���Ef��$&�ϰaQ�`۷�+�,=�a��(���
c�fpu���]�쯐3l�{���^ȑ�mv��ŝ(v>���RKŦԬTFr,R�fDj�������}��{N`4��r��{�`�7�b�'g��f���J�>6��aR��VJ#�agO��6�tb���PN�*�ۈ�hǌ,C�
*B�B,���n�4w&;�S�\�#.�`1��8�:*��Qs��� ��1�;��j�p�u��7�?�R�F�#L�"#�o��&�uY���u2�mHB�6?�l`\d��O��+��zj��8Sbc_
�}��DF)a�1IpzT�Tgm���THB�c�r����Rg$GP�|в����1�ԻM�-�T��ډo��i�I4b��'�(&�]�R�}_ �èF��l��?9P�H�2ƀ^>�� ���/�U�>*	��z��T9;��N8	�%ޕ�iZ	�9S���hB��P�\ۍ��*���-��0=����uBx���� 7"��T6��MN�k� �Ǟb%�>��ԪR,�]���v��@(��|'�����y	��s�u�N���q�SoK���d"��[��|NMM��K�W��v�5p�M��߭TC�r���n��'�hW�#��=���Qթ܄d�zb�{>z�KH��g˯�a�]°����*��p"��r*�%`Z����&Ѐ�N4��b)�y���nnwvd3F���.)�ܣ��^�hܑ�>��M<�	�:y� REYy��-���cQ�ͲDzcptn\H��$JJ1�z	)��[A���Q&��)S��.�r��O�]�$5\�_c�,�	6}��i����g�cfIp�*ӄl���_��;M�����H�p� 4�"r��՝�quc���u��㺖��QX�b�W�#'nr�����4ғI��g�)�A2ys]����I�� �d�P1D��7�AMQ��b:id  <{�����9���NI�w!X+�5�/1onϰ�0wv��DN���9$�|���\*dVL��܂3a�x5���Ď�� �ڽj�3n�~=�\�:�$���h��e�r���F��.�!�1�0tk�����F���1s+{9�nׅLB��p�R<��;���5�Ż��+�����!������px`�v�D�p��P�f��˨
�w���]6>y�(��4���xR�������S6'�B~����j��\�"�֫N��It0�irؽ$����̶�J�w�y������]D���)\�a[5y��Ѽ��t@^s����k'����+;�4����V58�y%��P.�n(�b�2���	L��!J�\�b~P��-����s�h����#Xl��Z��1��<�b,Ҹ~��6��z�,���8H�'_e6.�lw2�	�/F��yl��!�$�LU"Ж�:y��|Z�o�y�K�μ�,�;XY�;0)��2	z=����j��s��y�hh`��\v�7e���D}�|�ʵP��Q�~�mJz �^����|�RT��'G��#��r�6�0㽳��e
i���q��Y�D|hX����\�~�V�@J�:�y$j�֥�5�E���t�V����V)"uE�<����8��;���,��Q�K��J���u��O��Ӫ��V�1�T@�틾�S�V�84����lB�#���P���LdU�Χ���k���P����k!�ϼ���+ӏ+�"Q��e���B�@�m?Fc	J1�Rc�.yd.��-�%�fc���T�f��V(̾ؼ$=J���=U�����\�����m���j��m.�$ѫ�����/�����l "����E���s�����n�e#�y��^�; +ԗ$�Pf~{K��D��~�űn�=�a��\bNZG��r׸H�٧]xރ/�����Z�zhQ#j893-io��S�k��F~���:H�!D�=��o��>Q��|��v4V��<��>���?m4�?�2w��J����o��8[��@���=h�~@>��B�K���̗�˅��H~2�ж�)x+��qsG���,i�TH:-���.�'dat%�}�y��
��"5��d�c�W��3��~���?@�$�3AP���:�gi��Zx�e����&�Q�9P=3��Σ��@��b�,�O������*9PU��G�8�!��s��oK<)e�/8�[�fZ�Q�-��/83�����/fA�L#PN�qα�8f��(Wlb�# ���'��&�̱�\�D��֎��r�-��S����6�ҲYw�;���8�ΒG2r��QO��4��ʇ��}h_a�o�(�j��}vn>ןw yF�s�cϫ���Oe���4�u����8	�sSd���Ӓ��֪�S��l���uS�JW�
iI��#"|�A�:�/tUp�g ��=~Q�w&��آYmK����v�to�o����&���_#��~�lWf;j��1�Pҧ���Z�i�΂��g���=�xVW�z��]-���ɘ,��xȨV-�K�|B���=8#R�N�N�-�͖
�#ʗfZ�
��7�~D|�B>�.Z�l>�Э���pkZ��na�x�:FPs�GR���i������A��.*��c�������W��G&�'d3��D1>�q�qE�q�y��R��02��t�ȕgD�#C�n��}UjPɰ>(�#O*WB��#�*y�}t�>�����B�*`P���Ce/۷����<��Z�mV��϶I�ee�w��u����
yU�LT�=?����_�j�Y�(�7~ ňM���Q�Y`����mv�>H8��ɫ�������"����l�0�%m�!��=L��̚��ʍh;����$"��N�k�-�B�� �gJ������b���ɣ) #8̋}�참N((	�ا�U�w�"o�E�5씮vD�چ�y����-�oǤw��s�f���F���.���-���ض�0�6I����e���.q���_��A�&�ٿ�E�4[���R���p?����V۞�Ŀ�ph��1|l�Iz�p�����%l�w�ţ�;z�����"�{�%��Z=_q�c܉�q�f�Q��-����]3���=^��Ü����`Zv9��O���a��TaAgR%�jt�6��1��r�{I؃�?�����`��b��B��������>y�ּ���8Y,CUg���6�Mst>�f̱�wN�8�6Vĝ#@F,^M�*���B����"w�`7S��~&S`�A89�:~1�,!'��i���4,OT�S�p���؝�?|$!�LܖC�
��&��Y%%�u���c�6]���p"\�0�OrM+��z�O8�zBv=���a5�p�K�Ol8��O�H����BXb�W�k�3$��2|k������1��M�Js�o���ŀ�D��4�S�'+�D���Rz8�F�ޥU�u����9��*H�a�{h^�Ѳ ���J�1�b��Չ�/9NTԸO��	k�%��I��-m������h����Zۈ��*k���i(�K�d�}~u)�o� �uĞ���6H�����kʎ�/_�*��)�,E���th�!L�zyŌ��Y�l�������״��lI�GP������z���OM(� �N/��3�v�]�t�К��C�ܿ����n|묣O�����8�01��dz�d���b,tsz]S��j ����X�S�0�����Dp=�r��%;���|���N/�!�ƌ�4J���]w��F�Y�iB��>�"^Լ��G`�V��<��:��mR ba��Q�^��cL����x�p/8cHJ�;�U��2���L�2&{���8Ԁ����HOi�RZ��\7�K��:�6x?�if7��PG�(:#�**���l
&�_?��;H�� H�ۛ O�Q"����xa�q��W��23��.#�Sb�X�X��rq�'�����(�4X*3$!A�N+]RC��d���.��[:D8�7(o�LwIb�i] �G���W��ĭ��6I6��X���*ݮn*��02ڣ_���pk��W���ؗd�O������=�5\�ĩ,��{m�ژv�n�����WR�:�;�<:Ѐ��T����Z!�î0El���~F	>��l{T�� _���G����S<�C��a��n^���4˚c��{�e�� ��?q�kD���}Ц�¨%�X����]���Yۥ`OF�����ɮSQ]��5�~u񀼾�(;�|�W���1�凭4tKg�rS�%�f��񘕿������A�N�3����l�ܕ�5TZ����n��,^nrP����w6+V9ˇ8�)Vw?�������n#>ˡx��� L�[�JK|�bY_��?�=���s����� ����X�lZ,v����!۸^$6��9��í�I��c<�_���.�p�l�2�Ĥ�F��y�J�����$�Q"K�:T�]|�Вo,��Kה���8�X��0D�2�ŏ��~]�K����yn�5�Ե!h#��w��7��6^v�D���e���v�QZ)m�K�y��R�OW�T��GE�j#Ӻr6=�0���	�w
�)�LogY|Lh����Nk~ۇ@/z���HN/� ���Kt.�����u)}��E?$���7�b���a$�,Y\�f��F �J�1O0������K��1��\@lM׾��JV���ﺍ��!�|U�����j�L�|΢�y�H�����k�~�zz��t#��=����@ӊX"��?��/����ߺ��ImO	��&��)-�.,+��W
c�\*��m������\7$�U]�����RX��ʅP��GF��񘚏~��<��Ͽ�ϫ�G��rK��ke���l`�3��E�ر�R��u�Jn�z, .��ڝ5;b���ȁfY埤<&��(~����ɗ��C\}@�Z��r��j��/>��/ك*R��A���T�hl0�j��)ڹ(m��Fy'v�Fpu��$�X�ow�>,�|M�ԡ�V�#C�H�|�v�4#�2�0�Jݨ��@p9�B[�ˉ�E�hǓ:@Yf�B;�-�����b����X-���u�+x��*�GW�8�1T�!�����.��a�R}�����
*)*"��d�UXW�83�K2���`@��N���%���i�Hx@
>�������P�U���?�Y���~,�Wℋ�g���9^f|UBU �S��i|z�Jc<dx
/Ӎ.Vk�Z���Cf��J���b=����A�j�P��άWIf릮(0��>;x�.�v�Ԕ4�P\��������U&-�7� 7Ժ���ҍr�p,y����(2�&�)p�O����}C#�Юi(����xp�>2�� 4�}s��&��Ǿ9�TC�4�������m�.C���Ԓ����m���hߌrX�E�]
����ޜ��\�R���U������T S��~L�=�C4�]_6K Tק&��v�伴�(�����!8O�:Eݯklr�jY�}�+�h�U> ��ݓ�sv���)��Y�xq�wzZ��-�x��ӭ��qaV(?��}{���d#m�.��NŞ4�#R���fUAf��t�95iD7�tB�7�Z��<�EG�f�kU�����x��&P�D@R��D���ذܽ�.%r�6 ��Ҏ��4>W>��&Є_dn�ټ�qM>�Yuq�����K��m!:�2��tɀ�gߢ�C�!8��g!P��(�8*����]�y�@���h�)О��`�^�/V�g��.D<ܶS���I_<tee����`5�'k
Ts
L���?`���sj���(v6 �^��橵�»Q>+`�	x���v��8UJS�㝑v}���41R��l9�K� B!&Z=��̵5�������$]�A��U�(�
BA p��O��i݌����);(�8g8q���!N�g��a�p�Vߝ�� /��Ͼ�Dr��t�����%�����#�A�?�2b��y�x���5�+�q&�Q�#�Awe_hi��P�ю��&�c� �P[O6��R��K���U
'��B��0��S-�b��|��zb\���"�b���]��r
�c�=�{����ۊ!L�=:�ٞ#D�@��f�S���,��bi3��я��^~_t�������v4|�8��0T|0*R���jO�q���"��vI{Dpoʚ�B��``���b	��~I��dp�9	b>�,����E�GgE4)6��4ty(W�L�vN�f�C���c,y��*8X�B⸲�䀃w\��S�Ԣ�>L`��]88�P:����Z�"�:`�'�����p>���#%?�����L+���W&��Y��tu�&�~��?2}��\���Oԯ+�x�z ��8�����������,apf�pC=.�J��M�H�I�������N�F&$���|L���x�1w�sMz%�܊�f�:���4��'Ɨ���Ro1!�
����,���>����9�V�HT8g�v��^� :���e���4!���Pp�jToV���D	v۳%Tm&�� ٲ/����?������pۃ�x*Ɩy�$6�f�3���(u��$\� m麞�¡6�q��Qk*�{ǔ���m� !�,��(��&��|P�5�G��e��ȕ�}?����*�OA[�g��%d��^����yԚa�M�^�'����v�4Z��U��C�fh��hlnW�ެ�g:Y���3s�����8�d�D�b��tz8{@��ɯ WЋS^�ڋ1���pX<�r s�%����Gж�N*00��p�����Twl��F��ᄤ{���I�^�03��Sn��/<V:o��R��������bcG史��qp�!.Hݸ,J@�=�0�m���0l&v�{�߁5��i_�!O�\M5�\r�'�b�`6s�i����G:C1h?�*�3lE�_���;C�
�q,GH<f� j��"h ��S6�q�#߀ ���əG��,uX;n�ˍ>�'d3�����4Hj@���WA�CC]��n�������Ds�7ü3Gx�b��� �s1��?����[�~g�IqzrXaѦ�%�
n�'�0��X�zJF���2c�&u�d�s"�Ґ��5Z?�ĥ��	��s����7�: �R��:wG����Лzc��yL����!�u�0�>�����Fd
W��{o`��{���������<-�t��Y��M��)A-�o������V�����V�f���aI��@��c�]��6�������t�Km��h��Sl{�I�~Ptc���[�B�RI�Ɍ|k�B1�tfb�r�Z3�A��,�t���ٛ�	�BQ��A��ե�W?�5/3��2���SKQ^ia�9�ʸ2��+q
���{�V������ۺn����d�d��L�9Jƻ�b4�פz C��xs�Rr�;���McaX�&�Z��Fz���6����6���0O�%�~��_[�u.��l�R��?
�F��y"�O���?$('"Ʒd:/
6|��po�~eK�z��݀X�E&0_Y)2�0���Yi�������i?c�/�h��/ے�7�z9��D�.�� g��QyUm�';��(����2kT.HG��#�r�c�0Y��$�
_v��'K�Y<��h�C���`�~6�@�����,(��$�릦0tɉ���n)�M�E�+T�	������<V5,��Yh�A�_JH�=뭂�����啊�[1�$�@�ھ��VE���ة������ﶦ�����L�
�Ν	B?FX<1X��aC��=9�OV���)UNӅ"����c���-��6��m���	�C��˖$�.\��Rc�i�Jv��iHs�4f$s�`��[�٭�
���\��ۂ�ޚj���w���Z#&�ѱ������&:%������[Eh������/nȯ�{"ȕ��;6�0�?f4o�Z�S��~�� �$��מ�\���Z=�2r�����֧���%Ҝ�l��ɏh�]�j.�����cH-ȡ]�Ft��ޡ���%�s�No�2">�M|����<�V��E��˥17&4-&�2m��J���{a#ԙd[���s�h���@tT*B����en��A^:�:/k(�Z��`�x�&�MGҝ��`]T�(��-�2.���a*�}�0~�K)
�p�"�ޤd	h�Wr�3��a�R��@<tKiU�F�����i'�Jx�΃��U��l�P��������i��[�,�_�&ى��>9���U�"��n������%�P<���/n(hQYdZ9������e�!�ݰڥ��A��P�ԑΧVfFR(��Y�s����Ư"sB$a\'���v:PY^-o� �}�,���h��=��T���F2(2���"�j���}.�}�#(5�i�s�.>�2: �/�s�6ϡ0���M�܏�Q40�����r����R��и]�|~�������I7�'���@��
�Vș7��w��%��U��I�hv �q(~G[����CK1���w�v�tZ��2A�Î~���JS�j��l��j�S��(�Đ�X��oH�ĄM�&�s��x��>z���-l^��O�خ92V#�2٠�J�5#����N�/��C�M�YBfP���D����DRn<B4�SZa�
�F�܏�QkPqz�$��xU��P���R�y1�5�[�w�3.b6Ƒ�<��:V����W�6<&��d��4�z�>�a�q�����>�1���2��tYmgz��C����3�P?��(�m�*M�H��E8y2$8�H�!����U`��r�y,�/�޽���^<�����Ё}I��e R��k����
/�Lʂ�?��@��TjJ��(1U, �T������QPB�`!�8����vg۫8����~�����p��l�ڿ��4!��=��^�� ʃ��1!$���M��#!�BiN� +Ǖ�/���w#�g}g)vMN8���P'N��KbN>��#���x���t�
�D*��o�O�l�^��q#�T�.��m�?�T���	�<.�,z�l����Ee:S�����;��8&]z��q�[ �ӷHA�&KIĐ[�N'˼��&_m�g|�Sz�s֒�>��K�@ǭ�-�������6���&ڊ���=ł�ي����f�u�������3����=(^Y��m=��j%v/iL����׻xT�?uRަj*���1֟N�l{?(���8��Hr`���b�1��j�����Ԙ�>_~�r����s�b�g��)6�]Ft�����MN��x��Pd����,��|*�+�B��߄Yw�RS���4w�`b	�8S��:t%�����]���0
"�ٮ	5Sp��3��x?/���LRߠ�@#�&7UY�!�uc����aS�X�\�kO�z�+���z{U�8���al��ղ�a�0dp�N��E�B����Hs�P���<X,��!��$�o|��&���y1ҢM5 kܥ/�������(x4��'a����R�k���� ��k�ŝЄP9BXH�E�q��^O|� ��������Lؾt����.T
)�A�	�kB%	���3M��V}ʥ�b�,�!���~l*!R���A����*�ss�u���_h }鞥ɢ6�W6�~{kE|��(���2��[81,{�����_��4��ҭ��9M�b ~�X�|�&����;�b+�����\p��8����M�|���;3�(�v��#]�F{C��wV�n2.�����?�.G���5����d��b"�Azô�<�Ư�v�N\-��[wps��r��?%���2T��Q�N%�:�swԨ���OTw�o�F�uh��� �t�U^�Ĉ��fv��i:<)�l:�܋R��A�Z����N�cBD˲U�p�+�H���J����G��I/����&q#8�:�v�L�����bO_��\�n����@6n	�i@d��f�^H5��g*�P�l�f_u)�;>{����H�� ���"�e|�.+�q&����A���$(�	gX���˨+'�é��H�4�:�����ACY�]Ȥ�F���)tќD���7^*�B��bK�� Q�R�����Y]�I�+yX���� ��n��0��{�����f.:�ea1�d'����G rJ�5һ���>{�q�l�N�?�c�O�x�M6�:�����ж�w�J�񅌳�!:H�0EX2��F��"bz�{��?���0��k2�F�	<�,u��q����C�,�Q�Y��1?��!ѣ�G���a�Ia?l��}�[s��KO]���ϡ���V��"��ڛ�#ېS�H���|�~+��4�q��M�L�������t�}SrI�L�\"�g��H��}Me�����p�����\5
,��m�����^dp���ּ��T�+��Ї.��Vƞ��*#�!��nҰ�.���L���JA�b�椵*<�Q��s��^�"�3X��Z"Q�U~�l)�O�;6��D΋�������_ֶ�.i�bl(�?��QlF�8py}_L�Ir�$CĢ"A��:
Z^|G�ob1�K̀��=��X���0z�"2z���T������Md���vih��ۭo%7���� D.�����Ɏ�Q�p�m{�������HDk�TixfG{�
#�Sr쩨0�G?Ot
��w�GIYwJih)�w���~�J�@{H���`#>����M?<��tdSC��k')3��E�S�$���X����,�V�9��<��J��L�`j����A\��e��15�y@�l�����V���e
���!���V��5�Q�=L5*Θg��c������A�p!��*� =z����SӀF�"b2�?�����0����m���	���#�Ζ�,.���V�=c�ѿ����D��o�H$͛����uG�@9-�&j���Zp�E�ܲz����ԫ�;g�(�3��.5��d�)�;EC���ȡ3��n����M�P}�;Q0+��]�fy���%��~�9��1͒�_\��9Z�& rhW?�0�.��� ���t��_�h���j������C��<��Fos���:�RFq�oomnI>�D\|Ìn��~zV�D��������4HI�2��J�4{��r[oҞ[|Cp�λ]h=�@�b�B1`��@o�|z���ҵ#���+Wox\�����%GM���YT�O�Ȩ�.�mWa�)}N}V�/
 ��"�5�dD�W���3����J�@�K��$��`X�ˁ9ib�`xv�a���!�b�Pn���r 5�%��,7���(d��b9��U�>�0��_�� ��<��/	�yLg�Z�Y?�7����u�XD��^�}AP0P�΢�^f�wv(���tw�$cPƊ�A}�\�����|6-*5��6㈺��.�CHx8�bP���2��t��<�ȅ&����}�
�F��(�>��n�>�k ��Zs�r���Ϟ}����7�4ˊ]�돈�I�o��Y���n���Ԫ�������*�;g{
zW��T����z��GU����C� �2~B��7��ʔK6.�`vx$H� _�ܜ܎����o��%�`l��WjO?ق�;�ˊ%�+��� �xv�.�4x�pzP15-Gd��I��I"V	�Tf���#���$sN{�w�~����d�fK�љ��ܵ��gDmLB��XZ< ����F��L�kK��u|xєP�LiR���s�W=��.�v�����?�!�/W4�&�� d䄣�{N>���qV�]�AQ:��u�2�q�t?Q'g��C�筒��OP�)�(���*��HݴM7ym'���ϞS��`���Ӕl�/L" ��t�<R���>w�
�Ime�26����$�

�L��?�%�{��j�sA(�� kf�y��w�1Q�f_`�@1���v��}8˽����l��ֳ|�Ⱦlo��˃!�6�=}5������V�|��$�K4ϒ���BĢC �A�Jݰ�_2F�B��)��	8�� ����N9F�?���ߓ���x\�E?uD��W�jb�����'����~�!��������p��j�����<����7�fe^�C��ȝ���&�z+�v}[;5y�����\���e�Y��hс�M����|���z�|�z�KԆ:9�H�5�~@��Y���'��� �%�=����5�v]�f���>C�آ3�ȏ��^4���Y���1D�v*v!�`D%Œ��T�nHR���j]�l�����'{: �P`���`��b����w[�R���oH�>��͛F�B��}��g;e�6o�t�n4̂��N�"�G~D�Tj�,��*._B�^}�Zݢw���S��<��Ͼ`m"8nj�:�cq��r��eǘp!��F�d�`p�p��)��?��}��L��ݤ�~�&
Y6��u���Fc��U3<I\Pn�OCA+ʌ�z�.#8?�˶��;�Ű��a� py���@;���H.I���w{Ӗ���y�$3e�|<e9����1-ҫM�:�����u�g�Ս�4N�]'�����R%�/i6��/]3�����9<MmH����lZ^�� ��ē�A6�*���O�����T���	�A	,Q%��k��fɲ%�ʀ�T/�����yu{*|-�蚈>���I��Tu��!��X �0P����6Y^�9՝k`�-ǊTՖ��dԖo�,�T���e�2F���/���-�ݗҢ3�_�a?�ׅ4��]���3��C=� ��ŜM��
���S�ñ�vܕi���˸%C-۱��c�n�U�T���\v�)���A�Օxd�_b��z�*y�w4�V��Izd�A�ؘ |p�\6r�{%����m�7��N �A����e%B�[wb^�Fx3�N��k^�x��X����<D"�:e]R�<:��~��/Z@c=�B��3�p`UH[UJ6iz�昜���&���&lmP��t��� ��O�ۆ�_G\�����6i"iw�:����y�5d*|�!l���_v�;9[Ċ'�4H��W ���"^˼�	@+qad��V�����Ėd!�X��6��8�'ZtI�e]4����)2�#zA���]����>r��CO<�D�q77���=�Hb�*I +��4�7��X��4sNI��X��x��n;%0c�B���i�Ῑ��Ķ�d�u���� �5�=���.�좗�)Z�K�I�H�w:-�W�m���Ѣ��Ũ�g�,!u:�0��I�yF�I{�^@�qVC�s-�䁇�<c����A��K�f��GC���WC����\�w��H�\�@��C�ׄA�vy��T�]��4�
��1_����h����S��o�	�Y~�x�o���H[��B͈帘�t���r�wr����̢���Q��x���R�6�I���#��M�	5�DѨ����B^_� ���n��.�+�@���8V�b6�eb��Sn�-��W���k>L���J���b�K��t)��-s�����X���"�X��Z��0��N�n���+6�4���z���RB_Q̃.D_�lc��u��F蓁y���x�$^��"�Xq:���|F�)o�5KȦ̚��FXEG�0��2�g�oс����S�_���MhTx��O7&�g�DiҜ6�N�J�Q/��m6U�����I ��CT�9G�.#��rG 0�īZ�^
Uo���brY��h� W����~�ۛ@6��崆�tTޡ�wTTt�<����)���Ep���?e������,
�7���7x�J��{a3v�&�v��ϕ@
�1puV@=,
�~_�V��? t��
R�xE��\���T L�?EΓ�f����#��A���$���xH�_`Q�{�t"�����*����,m��r	6�����	�.�����c7a�@����~̪��$�8���o�c3D�����A+߂?N� zP��i�ϐ�۫��H���J��C)�����ׇE�W��I�F%bn�y01z�5;lǭ��]f������C����~�\���m�M�#\�f�Z3�yrC��k ����T�R��F�h��j$�N�(���^W��B(FjI��W�=��q�qwo��\>��|����rl�V��>�Y�襧��4c��2cĥJn����'
+�[w��)��h�7G@��hB�Q���S�����p�8ն�m�x�X��GG�� ��$T4�I�c׶.�oa�jN}	� 4U
�_�"��kd�ZWS��3�R5���@�C���<3Dͦ��i�;�x����eX��z�P)~�:L�����z�1,r0��\���OC9oM�Us�����U��j�<r�/��cG��Z�F
t���8����Q�9�eA��P�?�Ν�cf��(C;曏����a��e���>\]G;�����-��}�Qi�"?��}���!�k0�52���=v�Ƞ�l�s7y}�.u�,(k�<�i_>CE} e��s��gϗ�X�X�W���4f|q���ZF_��'�r���i{��X��](��6W�
�Fd��v��Ȋ��]Uw���~�U $��~=���2j؎0*KQKE����vS�[*�w�͎j�K����ql�Ɔj�J邼�L�af�Ɗ������ՠ�lx�c�zˇ�-"�Ʉ���*V3+���˰���#���zNV�����a���fF���g�j�D��B*��Z���ʄ�7+�kF�O��f+x��!P� �R��S�ᡡ�?հ�:b.�;3�GՈ�i��2��W�a&a�id�&��/3>��q�
B���zU��B;2z��tzig���C�����^�P��<(8*C�ݏu�y�JL�~���c���: `<<�ӯ�}/ǅ.�sG�<�����lƳ4Ip5�e���)�C��I
匾L@�	?1�voAj gT(��j 1�s�R��Qƪ�`Wb��B-v�8����4�r��֎P`�l
(���.!7��=8����?�y���W $���p����B� ����e�`�����k)���88�ܶ�pN���Ce������2��Mt쀯�DC���e�0������̢�������sL�J����E�FTآ�^��il��Ise�����!��܅�&�O�1��[V�&�>������^c�x	��4�����퓴|�O[z��N�U h������u�y�#�tσ��i�30�y(�2��so���N����@��c�{��~-��I�)��mQivސ�#�f=\�$G�Ѣ���Y���}atlf�&��;]���{��R��k�*G�<�g���@e�fp��K�ox允��(��a�
-���8"p,Ś����	���S4>��50��O/RZn߱
C��z��Z=NR�E_�!�^5�g.�s�����1�:�,� �Ĉt�lw�7ZmgCDl�}��|Zu�y~�A�s<_O�tX�hjZw	�(�c�����/��AC}�������f����Q�(W0F�S�7��Y&�B����$(�ݕ���Y�FĠ Em���,���Ķ�6F�)(&�M�������T�O�c"N��<��]��5H�����v0P��G�O�h�B�|����3ԣ�ܕD��34~��1p�i�n! �`jPC��j	_��O���N�"nz�HM.��63�D�|!�(ȼ�@*N{����o����8��ݪ�6�}��AH�9g~䐧tJ1|f������'�˅㔬�]z�➨�@��狵�?"=W�GP�r�(˲ME]%{"�<b/��o.���7��l��{�Zp�O��������DB�e���7ƌ�<������n��-�_ �#*D�Q����[���<���5����~� VC�8�	8b��s���t6�j�0���9�M�5�i�i�ހu���-�̤pm�%=w/�����şq/{&����DC���q��'RU�3�R��2 X���T�����g��b�� ���R֓��kdvG����)�|R�/ɽ�&Lo�V�0��sy<��:�߬�!�Qg��>���-�Z�g}�yC���_sK�|��X��S�[�T:.��lC�a]��/�7�w`��-5P�S��_ػ�Q��&UdM�o-5�?n��;`�/ۅ}9��E/QD֍�	��#��-��#�я�2/P����TO������o��d��?�k�d-\5�6�	�\-��Y*�d�ۊl�Ԣ��]��H���Y�n�_����nVFϥu�x�s&�-���2u���V/мw�nA��Sr5�
��!�ȝyIi9
����@z5,�EC#�:�a�ov�ȃ�^���.ZY�Ź��"}�}?8���kZS��g�ufͯ�o��R�E#�"����4�b��=��|3[F��oRf�t����mhF �J�IG
h�|��!@p6����G��@N�7>seIR?���!�v&�k#p�$W�M�TQ7����ɦ�0%�_ѭ�\#�4!��!@u}
4�������>�#C0��U\-�B:�!W��`]�kTf������]��q���Y�׆��XD/���n���8��;0�r.^�Y,��܉E<)!�h��d�tq�r����/�T�	vAvU�	>ܓ�Fl<�3l���O���k������z[�7�>؏e#��P�
�os3����9�(����GM�݄�����e��֦$H����.�(��*�&����S�ţ��$e�r�*�(R79j]6ƅ�?�dg��Z\�#(W��p��G��N�L"G�mN�+?5	�D����DO��<Y�P�7YpLL����=~�R����Ɨ� ����^��n�&�jj���2��3���+*�Ch�q.׍gr �����M���2xUX�E`�8ω����'�l "�(%e�0�e4�}��Zwk�;E7�������˟p�����y��(�EEZ�n���?lу�e���AE��ZJ��W��1�מ8=N��<�B���S2 Y���F�9�%�Hc��o��5��\ƁOSf/�F��[\̧\ʴ�/���| ���?��h[l�	�T�[%a.����cl��75��v�w|h��6�{��AY�K�ª� }5��L�����f�?�ߏj���'F���f��s���ș=�?�رn�I=a۫�����霗���H�b��1���e?���vNu���{��sh.�2o�u�:���5���* v�P[T�h�;*J�FТ.�q�_��҉H�gKԯ���H[�{������-�bH4����=*N���5���k>b�Bo/�Rn�`!w,�#��ٞ*v���>pN<l���Y@���q
��awQ��|��X�N?���Q�ld�Z���(q)��'C(�o|�ީ0L?Ȣ�Q�rZ�-�#E���O��+#�,G���Ep ������}08Zf�ك��+�ð �6}���Qo	S'�%C���V�+ڜ4X{^�wLРr�A�}���Jdq��B�Ϥ!>m�gخ���T����r�2����,����.��km�EZ2�X�?C��>T�Gt�U�����Z_4�ӫ;�T���u!U�Gip�L��C��S��S��!
,/�0
Tf���3�^C�Q�$�Ť�^��!9]�f`ay�ȳkrMX�6Q.��� �1�F�j���xߖ��0�Q�:��澀��MN2�~P��z����2Ԁ�-X�<��)��R5]b��C| #���������	æe��U��0��b�5�|��tqK�"�9S�]�¯2�D��|�^42@���GK�J�����aX|�N�-�-0��q&CwvQ��^���2@�[�l�Y��c�Ϡd�&��uS�j��(&�GQ؋p��F|�c!|��P]���-�tf�v=pN$~Zy�p���4��#>1a����P���_�*JvY���,C+���������[ǽOX�y�ZZuXXp����:bU2����yxԿf㉀E��.�я�k��M_���Ys��T�\{�I�|��.�J�o��@��1_��݈bg)��R{t+� ���B�Ќ�fU�!�\��3ޭ�;y7q��a�BÀ�U�N+ ��'_�&���/*��R�n��'wG}T�C����h<8�O]"�P/�#�4p��E2����	܋��?d<Rc��*Δ�㭔Ζe�e���"	sğNׯ���lZ�|�$���v�9�|{oD�����u�t�i�瑊#���sh���5�0��p����J������X	��,�w���ͽ�Jŝd+Q� ���B�����6�nV��{J~��OJHz����\K���A��k7��G-�����-1�()�4q�o�2�����|I1D6�� �۴��~&_���q���Q�C�����K.~Lڠj�<3����(8/�5GX���h�K�����_��8\C"�%��f�XW�f}E�;�P{{IԹ`��N���%ݓ~�lI�}#=��gW�<���&s��u�jĀ.�c��='Y�-�ڡ�i���Q�U��9߼٦�.�d�"ܱ5�X�G7}���fF:�{d��k#�)����t*��{��*Ĵ��Qf��K���x%�J�:.���a��>�H�H8b'U:��O=��V�Γ�p�&u��wTR�}��JO���A�ȍ��R���_5�^G�/gnK��+�P�z��,&��Q�t�+�wyg���l��Q���V��ţA4���fOt��g�AVI��������/�X�A�����O>��ծ��_�'_Γ�o�!Z��id�Dng( ]+�^����`��mШ~,D�����6��/(f�SM.u��SA�1@�lRcb[���>ߺ�t��\4t�[�p�FYP�d���y�J�;?Q3���Ճ��s[=�Aԩ��!@��`�ĩ13jI��܏6v��e5n�=�Mn�%6s���(a�h����{�W���+(����"�6��T���HP��g��z��s�1�M�[|��dw�%*���]�N��R�'���f�"}f ��
�겁���]e*�"Ծ/�|_.���7!9�*�cꚏO�߯��r�F�(DUe��97�<��Q�3ZW�
u��<��c-MD�P����֛���|WH�Nm)�t_�kyV�@��IwMb�4r����lv��eo�xT����ϩDS� ���`���Qp�҈=�Ni����`�����4�Y�낊���M�RF��3�#�rOΚ��^��N���OW ٠IR3�����d�u�� ��DD�ͼ)x�oب�fC���
0�}�y|_!:�U�Π6Q�>�2,�d(�*g��xy�����6�K	<ʘ��S��Tz���˅롤7;_�7�`ơu7�S.�<���ȥ�Ţd�Tq-urn���`�nf�S�,�U�Q���I���c��-�Mq��h��r���8Q��2��͎��<��/ok������5	��Ikm<�Yj�S��G��;��(�U�����ǩ��XnU�@���g��&؄�8Fd2��b��>��PnEn��S���X�R�θ����iyq���N@�l	^*�̅J�z��֯M���z-�?0�Z�^A�*�"��D�`��ŜZ��-gZׯf� o��	���E"]�,�K�4�Ѩ�}�8|s�+��E�o�u�t�"��G9 ��I�q�
S��|�`�!�����G~+րmq7~z�I^A*��5"�A��#���$�fH֔���2 ���L9	��0e����#�E����uY_4�{����>�zj03L�U�/�I3!AN��<2k�-��:W��Vϱ5��Q�l����X�fA�(���<�ǜ6��;p����� m�K�8�ɼC)a|�h��&����r-���É��v�E�Uʳ>3���q�s����O��
>�Ջ9�g�M.a>o�##��P��o���\G�9ҏ"�2������;o�ƈ�e��3�d�����hB*ܵ{��Eh��$G�T 4e��*@P7yi6ma?4e���c��W���S�ҥ�Lb�Fm��?uAD �\��.��|ӎRi?�w�4L�v����ޒn@�TĦ'����~.^���fE�j�ƒ�2���se��z��IĸP���~� �~��&�����x�LE�(���*YGg�: b��%��C�񽌗Z�J_;��P�EF��l����*=)��'(�|Z�K����ls1��մ�a՚����z_��8}�*�_kSB24ɴ�1Y�yF	x% ��&�o�WR��������SV��҆$ [���\
�^o�_�S�L .��?Xz�h��S	��[e�<�˭��lǴ�5�s'v�Nh!��Q"��ޒJY$���MA�%hs5���\��X�^�Ю�_�GI�*��'�DJԦ�Xs�D��=g6�.A�a��������FC�\��o�q�d����!*�v��B�?���Sby.�	���j%:ӕH�uv1��hvB[�[� ��{Y��R]7��-�qG'�&�;HD���v��ʝ%��޻B�PȰ�m/�b�C����*��s6����b'��ooE^n�ǜwl����*��ޏ~w�<���ۙh�1A��ow�'�|�v�ɎuC��'Qʛ��q���')F�pgG��3����[?*�Q)�ΖV��#�5ڢ���+�2D,���ޅO[�D���8l7�ǚ8������+X%�`-6}���<��w��GF�H8�ԏ]�ςʡ��)A~w��l=s�]�����a\���&�7�]�m/�`zz��2���哤!��C��%��`l@�zoy�ٻ�1r]]p�~�'
1z�Z�I�ۑ�iH~8�]��	F�x�@��n��H��ĥ�
�2U�x�єmF9!?+e�XfxVw�Y�����A�g{���/v��mb<���>m�<��5���fg���L2+I���B�$Ȥۦ)Fm��62�	?��>`G߉~Ȫ"X��_�/~N
����2w,��d��t�(K����g{���?)��n:����,z��:4Rk��ݶ�ț�n��Yj����Q��U6I%x����U59$F4!�C�����3c5�¢�S���j\�K�/Z�n�ˢM8�]���y�h��pZ8$�j����T�*|J�P +��>�7��56�Ol(�IS.	��H����	R��D�`i|��VeQ]5vR}x��^��G���<dc3ʭ���k��Ol��MT*ۘd0�ڽO��x�d�zRZk���˽��|^�Ei�,�t��x~ٝ�
`��i�����x��=�E|n�
�je"�nC~l���!��?��7=���?����b�,.�M�߰�Q�$���q@����L��a��'�,8KU�@�������������j���>�ۉ��w�J�Jp�6�O��
Q����k{NR�DDb�=� �/�
�2q����X��%������ޭ�"���A�M�m`�ri�����%:�ۺ=���!r22<ܞ�~�N�]O2�:+C���L�(� ��n��"������'��K(���a��m""3�Y�9u�&xۈ��~!4O?��aB����73"k��Σ�;�C�<��*-�Ӌ/� bG��HG/��u8;��r������yL�~���Vi�]H�BImY�i���n9�w��f�B�<��6p��po�ð#榝�x�p���Z^��zt�S7���\�����@G�\�'AW倥J�ɐ�[�����6ݢ�����*�mAT4V���״=���� ��C�[�U���ݤ^�V>��;�@h�"�B�����Q������(�qJ���^�G9�}y�l������յ��B�ڭ���
JF��mlg}Dq�B���O�+N�� W���}�7
R�[o���I-�)VLd�A���]W��C\C:��
��Ş�1��o�f�kd^v	.���J���Y�E1m�1�	�v��wѡ2�W����h�n����f���6�������O0�k�B���f]�\g ���^ٸ&b���=��%p�	AI}r���S.��e��Qdŷ�8������_�@춋r�.�>��uH�#�+H�K�#����5aęJ�.�OPV��[XZ�Wb����q���^\��=N}]&QM�XTU��V+�؃�kP%%�ã?s|B
t��Z&�C�]e8Z)�W)	�-p!�Қsݡ ��:-�ɲ��h�fM�� �C�KB쥾�l�&�q7�J�`&|�^O	MO�^<Y-���^�'�]��j_�8;x?W�w�>�^�u4k*U��x'X�,`��y��ʸVi�i���kd4�h�٦� ������ю����@-�xLvF{88�?nR�
)�� ܃~9�Ɣs-�%�7Ҩ���8��,�����.˵`�g-v� ��y����#_�
okIz(�0ٝX�B���#�AV���Iz�u���Nv�X�����K~�BT�����T0Bz�\8���0Se�a0;������� �gi�>!*�xQ�t�A�$.ϕ�$	���W��i݋m��d;�ʺ섃C�H�D������m ��4�'���PL�?�wFC��@�� V��F�TI����^u�P:Su�!���xYAtg��7|��`��0�`YD�ث��\���5��xא���"��ۊ�5}�[S���(�%���ڿt�<I8Fn�����<�04\1!�߹?�0�u�v^r��a2Ѳ�����n�)"��٫.� L�^/CiC�pB���$���Y]//�!�@0Z3K���w��8�T{���B������iJ�Si���	K�_��h�x����:i��H�<W��e��c��:����V*u��^."��Kp��A���E��~�"�/-��M��Ub�^$$sC��pw▏��x��Yr��֖�0��y���y�v�(���Ɯ��N]�(��J�=����@�c�$��ܮGJp�5W���V�JN_����Z��j�w�!�$��h�J��l�B����_y�d�Ћ����b�9f����l(}%9����C���*��`'/5l9-R~���#�Ŋ�N�wR<�d��<0��40ؤ����~ �y��
x��}~�e�t$$�(�P._�l ^d0E%M5�)���z�PR[Ƥ���h�X��́r�ʏ8�]� H��>z;nI߭�o��(+ݻ�Խ]m�Zr!��4{�.,�d��XM��3	�b��M��*y�uf���Ek.1���\��#�9e�s�2 �a|{���|�)�.�Үd��@B�y_�#�7�q)��{��. �-͗/��R�U$�&��9
���|���#4y���P��uġUG�5p�'4�k&U/?Bΰ��?�G�~���=���c<~�]��m/��L4%�ف'���}��	q�"�t}<'"L���Ωl��I�
���;��ټ	��N����mZ���9 -�X�ٖ��5{d�ިO�{Ǫfb�>b���:�
^�hj|j50�����	S�3����&yn]���1(�7�JN+Fn3�$�̂��Z��z��N��&��U�Jb}��� \����Q�]��C��C;���ɜ�q��Z�q(� q2����ĠI���6�V���ս�_x��q��̶N�dC�|����KC)�L��i������F"�G1/��X����c*�K�� Ј
����\8�%�mfFP&X,�}�2��e�I����莓�ct%rK,���R7�s��Q�S�t�۲Ƀ�I���dc4�o�NB-`���~nQb�wQ�-1�.���;.;��R�����۞\}V2�fa�X�plu٢qN���{*��b��s��5H�f�5K���x����ol/�� �a8�_�]/}8xZ�P� �ڍT���.���~�v��R�P���:a1�^�6D?�/BSR$�_
��^��Bg�ci��0�Ioh�,��Sˆ=t�?�I@��[M��n�=�&���C��"���A؝y��[
�j7|6Ɋ�{2���/s��j{��wDׇv9���A� ��2Ϩw��eD'=��u�,�m���v�P��c��/g��!�Y�y�[ьג1�J�������g��<GR��Y����B*�+򘤪���3�%5474��62T����K��1}�@�I��Y��3�Z����*D��f_�N
�{@mAe̜Ҁu�1� �b`�{����sO��H6����������_hT�G��:f�P�%���K�Ձ�������i�S쩆�9C�vx���Z�&����^Y��@�P��P3e;N�P��`q�)��e1ߓa����q�w���MV"N��3gף`���;�����I�[�FH �sI��>�|uu�%���7h�����D��::0˙���^��<u�<:�7�G#VSF��3Ov��"����gY���;M���j\D�}�$�O�,sT`(ѡ�Z�� ��)X�D�?��\Vi%�� ��ͤ� �y�����)1�n��9�@�5z�QfѰ�'�m���'$a�v�K絒;���Rb�#���U@��f�`�_�\aY5��}�cL>��j9{�KI?$݋�ע
�ï���vax���Z8a�j��!��8W|gy�z	ě���h����9�	��tHa||��.�RZd0Ľfhiy�mV1�5�%CU~۩F�d\G��E+c�+Z�rk�ؙl�H�1ٱX\�0�WO���x��Ww�Zks����=½� �|�JE��a�1��x{�N��&
�i�i~���dƳI[�E�;2
�rªyk�$	땠�[�B�7��|�\`߃_@A,�r?M� 6V�%$Z�q�%�1T��ȭ��9o,���=���S�}�1
���v$瓧��)\>l���O'oJ��������0Y}�d�Sk�˘aE�������b�z�Ӕ2�X2�Y%�N\�c�[���sq��
2jUmr)��::���|��Dr�0�9u�~��c��0�.��:�ǟh�L��q}���Q��l�/�5�#*���r_a�"����IL9r��&WP ��[��O�`�a_�'�N83h���L�;}.<����"�m �ź�H�9{���;&�o���\�dj�L\��!>V&
H
ZymV���)9�-��C9��uc��ډ��� կ�M �[( p���c��hG����S�����6V�j%�x=���I�A4�M�"�wɭ�I�I;�����َFt�m~�V�'�Tu_��y�Ԥ��XG-��X��M�?VId;���h!e���+8Q�D�'��(�\�_���S�}���H���yb[ղ�Bi���L�
'��곩}a�B�yOxjaN�W-qlغ�
/�o�!�M��ݗd��i�=�W2U\�X��玑�B@91�n7�#�-d�	+�����c�L�Q�"�f]�C1��vc�.;4�Tu1 F6g����y��	��z�#��h��{��K�]����/�{&۝�Y��=8���n�	~�rz��S�=j�.jݪ��?ժ��Q{�n��@)v9rj��׻\��#IA̨����[�����#�hP����x��Zn�K�R��q��>^���=��&.��0���¨ޕs�k����v�sujt*u�&��� �8wbWą���d�!�R�sz!��˭`Ŧ�<��DM���ݰH��C�������qt9��=�Ż۲Ml�����w���8�' wl���0�?ԏd췰����4�E�U�['�H�,���y�~��&��'��(u(4Z�b٣��zt�9�Z�������F8�LӜ��R��Sۂ��������a�s����T�ȿN�Y�ak��q����`J�I-�A�Q뵖�+�O{��g\hF�z�9W��F�BqH#|����FzS:���U㊏At�VYtB1�*�\��TM���]�,�W���-�,��d���a��¬ D�iz�*SƜ�x�A�;.l�X����*�W�7i��^�Jp);����sGC\D�_���Ϯ��%��	l'IcP����C���8�����T�G��f�^2��P��su�j��n�A��h��[����7H{����5V8�Y���B�x�]���HU�W�R�[�[W�%H��w¡�yn�Id�$�(��E��`������	֖�k]u湀^�n��:�ϊ��A��ˡ�"��J���v�=|X^{�C�9�p_�(��Ӱ�`p�
�؊$�x�Bupv(>��iic,������-vE�bg
�LG���t��,�t#��!	�7_�>��ՃDe,4NM���$�i@q"��֘���
��sn,dh�bDm��۝��І����8�Y�n��>Q�O��RJԁ�Ә��ԕ��i\�k�F_��@��)L����0k��YH�X��;%��w���`a �X�4�������r�3�џ�:��_��[��rԾX��6~􋄇�0���z:����ML��V ȔoQ��D���ۻ���/������a5�b"ĮȔa�	9�'B&�@M�0k�`g�Oa��a�3^�33҃���s;B��<l���5nӭ3- �ϙ��IH)XS�4��;�w��U���iC�L�ofK6VH�-6m{<��D�A9F��H��?DZIC��n	��]6���w� �Jp!��hb��a���HS����>t�Y�=�x��T�A9@��V���U��.q��;.���m�q�V��j�����I���ݛ�6G}ߣ�[������V +�;.�hQ�	��v���y�Q�ϣ��(��W�d*�iK�}��ʾ-/��s=��P�B.�4�\�<
,^�돀�}�	xBy�qO�0kN%GW����G
4cpo�&u"$��|Zd~<��-)�W���\��ѩ�D����1 ���[�d@3	P����(:ձ��'�m�'1_hMvH��� �y��di���O�D�N:��X�������^˰�"��]�>�B�����&��L�
=�xF����	���r;�SPM�s���C���k���\�3��@���roq��`�C�׮�#.^5�-J���쨿 ���;�)�/PxB�����ZS!��nq�%(^��=��&37ևzz���@��z��k20^��
�sލ�t���&��?8�UW�᐀=�!�;�s?/��0tDū ���
3M�j��!À-�R��S�Q�qٔJ�BVs��{�M�b��������'�n3�l���-
?y-H��� 7
4M='U�C'�5+,J�y����x�E����%�4�=���V%�?V����֎�l��b_��XF{i�!_R�}��G\;�%B�����sO���D�3�K�����X�ې�Z`�ӯ-�op�BC����R�4j���'���Kz����? 7BvN�#!z#�^5�z8>}��+�ztƏ*k���B66�Z�T���B�;�ܵ��R�e��K�8e��2 �[�iH��*8E��Vc�A-+�.1���qo���3W��i?���/�O;�?�
C!� D,�>�ͩ;ۏ@��x�'.j�P.�_���bCR��ȝR����GTk7�Kt^
P��u��C�3`~A;��ĝ�1�^|�^�.+�W�~�����uxy�4��,��!�����[�N��SL%?,��<+�����Ir��)*�5�E���>�C����VuKХ^��5��[��C����P"�="�j@��'L^��C@R�p��7������1Y�Y��ü0��M���ż�������i�W��Ew�5ZXJM�)�\��-W�󱙲�	G1J=�RWBSiV�	_��৤P���wb%�$�I���lK������_&(yd������-��a9�,l���l�iF>��c-��I�L����'���9Z��~�	_�d���H$P8��J��Y̫`�O���r
 E"��Cs%-��.�ey.Q$����9].,� �L�E2C���b�2z��\[�����d�����9�x��B��
ĽHF�~z(b~�:C��i+���*���g�<���{ӑQi�X�gU�`��bW��\�_y��Rf��pE���.�H��d����h�s?� �K�{M�g|��l.�1�]@o��_�>���<
).Z{6h� 	�0̈́s����UQ��^6H�Jyz������y9(A�U<�g�Ut����'�P�&,9{/세�T���,G�^��GU���ғ<zN�]�zv/IFq4rl��!��
�	�?��A��<�G�_!�Vi��h������|3�	5�Nٽ��^�Z�_���y����{�r{�K˨|���w����y��h��5 F��lڨ�FN�� t��9k�{/l�9E����6J�+�~��Q�h��7{�xO���(�=� ��JO�¯;�\�u����9���Pf����]���
�G�/(�S�qK��2�5��;`5I���6x���^��G_��qʴ���dC�4���<K�L�+��~��aKs�ݢ/�qtX#���p��K��{�Մ��E�\�ף%���f)�X��L}�r���QI���I���N%��V�l"��#6�$pp���T��W�
�&d��Bؾc�i{�-mEt�+j(�.Q�ȵ�����h8R�f��Sf���&�	k�}��fN�������X��ϒ���*	�i)5����f�dKBV�x�D��<�_�
�,aE�ɳ
B%8d��GHčP�����Ε���h$�i�R\�s�L�a�k��0�\��R�(�_wm�^��~g003���6n����,��]�Sɒt��gE.�l�S���~�;��A��'�v't��A,Zrƃ��[r�I��/f�AE�Æ��0]p�eP�S���J���b����D��FB(b�Qɉ:��àb�mNY,����ƣ�6�yh(�!�M����P�3'���3c�
�����GǞ����4>����P�-B��b������3u��>L��]��Γ�ԫj�!��`,�D���jKR7��M���n|2�MpV6�JD�>�թ*=��?�{<V��1�/��^���6),�S�H��g��ѐ)��1>v���ѵ��M���n4]|���T��Wi �L�"?A���=H��&�t�]'�>"�	/6�.b�X7�J�,Ȥ��DiO}=�����HXD���eb�*7�:�<��Љu1�Ȍ4�a���eՓD9�9�d}q�]Pg�~0Ǟ�f�������6V���A�bnG��u[C�'���ǃ����O�uϫ���`�)�b�o����p�oM=������hš�Z�'��v�2Y�}��3��O��R��3u���4�1���Z�=Kz�V�9�d�@ �\RX��e��dxO�������>��1ç�h����yo0]��y>�;:🿬�Q)�>��������wg?H~yE�r���KK����S�PT|�[ ���#t���7�9`ZJ���S�m�������%d�U-7n�n��r`I���������Q�����H��k-�Q����<�������
V�;��z��CQ5�����Ԙk�D)�
(5��1͕o�GY�_��)iዃd��Q�Xӹ].,�p x���n���g�!�z��&ڦ��z�627���X9��R��n�b�S4��Ej�м(�}i�}��D���o�Ɇ��9�*M���A�i&.&��R�g���0W��Vi�	R�D��;6lźc��C��D�y��)v�d�3\�n'C��P���/A�CGޙ�2Ε�TT@�`�K^,~�PѺ�u�q��(�tA����N�\�
��C�o��������Sx"~���mϖ!��[
M��#%���1�y�s�IO%t���nѪ=��OI�Þ�V�o���)u���^*x^�X�5щ�Ǌ��
�" ��_)��7��^Fp�C��p����v���rzY�"ѫx� 0��7������+1��~�Y�p��݊E'JB֩�b���'�~�QJR�{W���VH �_�/[�<~��$w7��$���,j�l �'���*_ȴd�(F�2`���:s9������lJ����X�3��(��s '�O9ϸ,~�/�EM�Lʇ:W�F���M�5���F����{b ����ǒ<�_�e�Π$�x0�@�.A�� ���E�Lɲ���QOz�[w��{���أ���,�����H��z]�)��[�g}�+���������;�t$����8�X������bl���6'yOUf�%�EM��.1}��9�������,�s�Ք��h�{B�(|t�F.7D�w�@��_�G��Yh�)mЕ{+U{ �W�͹qo�Y}�U�N�s�K�����&��+�y�x��ظ|��0U���}~'VF&��/�E���8��GX-Q���<���R</)~]��K/>��4Gy�INh����	���V�5<I��s��K�ѭ+���3��Q�	�N��DZ����D�:xЖ��
{�)b��mǌ{��`��a�D��hL2�55�L�A�V����`���ٕ�tI�.5>�d�zJ<¦+�f��Ʋ���h��-�!�E�˗2�h��J��x���\�	N�3�����ť���w�f�mm;�|Ao(�E�q�L2��פ�}I�)6m�"z����7c_ړ�q?�P�0�YC�7U�q rK�4�Lq.���s��6G�oT^/���XسK�ŋ�K�{G�jL/�  �\��4%!�f(�pXN��}����]Ik���iԓ��i%\�~,k�%lG����E�2Go��3t�����my �I_�
��|��&!�����@�����͐�7k�I�k̎WFR�7a�� �#�<�$D1$���ջJ��r�W6�02$�Z�#�i6�� �u�9B4�B��|Ľ>��~0 H�U	��l|!����VPk��c��8�ʮ �~��ξR����X1H�uş�)ѐ��q;��
��1_�v�X3x�v�v)��h�z$�A��rZ�����9�Ybv��sU�e]>iD��s.� tB�Q����y��"�F�Q��&�>e}~#�FPp��o�Q�)��9?�D�?�4�U�Gל��5eb�˦��O��lk��e�*�Fĉt���@-��A2e���*E��7FЄ6s��?� ��!��hWҿzy�����*L/jYm��?�#�D����0��i�2ڤ�LY���>ޟ6Ƚ�D�t�����E^L���3#�j^��?G�� �T�X��p�:���Z��3- �٩��h�� ��xB�|E�!��3�ͷ٫�m/ /�H%�S��B��jm�ZA�;r�����/�c�}g���+ȧ�ģ(~�$Z\���	�l�m�����N�/��2����y�d�a8j��좝B_]Z�`��Yz��F!?�%���Po��Z�{@���dS#q���iD[�Χ\� ����@ÿ �Q~?�]�hh4`	Xo[r`~���B�8jbl��%5}b�vAh�f����S����Y����72�֢5�)��\C%u,m��8�̲@�w��'sO��3d�s����k=� �%���	JahiQ��j��i�W���]�D��V��Y���O2v�oR�,Ȩ��D�.>���$:@�Â׽Ľ$�v�3�[���y��n�Яd?q�W4�3��H�#;��e�ܒ������g�|s��\�b����&*۠�#���� bT�o<v�n0�wy~G���?*s`�k0g<9d�ƿ���ރ�pw�|6|pm���A��QPQW�0$�N��RY)�|t$��\���6�$?��Q�2��#R�P��[�+�,4����K�1-����1��8g
��0�g+e���;�}Å<u��X�	F;�C8�v�]g��ʮ>1)��Β�,�s�'�+� ʎU��-<֤�7�z5`�A����g��L^���C�%�L��́�߇2����1��p䃹���z._�������~EA�][>/F0�-�����8�uFF��;�
)�����>F��I+R�|X�s�w��C��ŒAE��ԙܱ��)�}_�mmuî�:�����c-m28 ّ��n�qv ۓ�7m(KW299?�� >��G����W��i�?_�D+� Z�{�T,��u��JG�i�L��������!�!�⨮�T������=�O���z�=Ԓָ�!�J�f����@��rśQ��:[�p�ʮ�T�������m�N�&6���W����(KM�Qv�^���cX0?mL�@-ЂL�1���=ybewC�&cՕ|�Sl[�"��ݕ��w�0f�bEN���t���~N�{D���0ȯ����u*�;?@�����J������a���N8�-����%�w�?I�ִ�Ϊ�+[`hg��H�cH��d7#=m���q�(��JG�<p-�X�ހc�-���=ƵATtޙM=���~�վp;ŕ�K^���aa� �����W�=sǃ����]��C���ʐ��/�F�ܮB�{�l^$;1E��P�ܒj��i	ʇ�����l�����$�x�d퓶Y�ו��E~���v���k�6����v"BN)��Qy��m �~@�ecS������2�ؤ�y"	ˊ�#P璐-i�6��M�����ؚ�9��'mjtM��g�W2�(�0���vjؠHwA�"v�����j �X�2L�i�Ր�D��W���ǌjc���-��X �@�Ѭ�B�_Y�{U�I����1iO�b	�����Q�Go��Yqe���pS+慎�:��3˪$4a���9�3�q��m�Ж@�G��v03��j�uǼ���D�A#��Ng		@j�Ue��ҽ�@1�@њ߂�{�;�~)��B�X���5�z`�N9h1mk�w��m6���*K%P��	{�+9n��`��s9���x-��7x��v��[̡�ݴӆ�ve�(�N�k��9&�����.�^�������Μ*ѮN�m�3�}:`fTP��Ш㎽I;�w��F� t{�S��7�juh���Y憨�(���l:wƙĠ������.u���:��G }�F���O������x�gv���츳�TL\�}'xXO0��T=��C���b�)�?ꜫA\S��½��]�ḱ�T�����n))̻�nT���=�zc?�R����}�D���3Ǽ�������W��v��NEU�Q��W��zV�.Y�5~q������j���KfM]�Hq2�g�x��
^�6���8>T^jST���|$���Ę�T哊��)T5�c6�	7)�H~$���ښR���ĺ��i
RV?sY5����ǉ�ˑ!uZ�Vv�c�g��-�k��l�_~��uu�'0q��O�Չx⻚��k��x��ᆽ:@)|��EC����F�xx����۟
:sai��I���f7�EV�
"cN���ztF�٠�fҙ�7׋��-~����,�b�MpY���$��qq�jl�N�o�_8�A�@,�����9����؝�a�Jt�����>���LqFJLo����������k0��Y��WQ����n��PK����X��%V|U��z��q���	C���y�rC�t���:Mf�׌A�Ӟ�rL�j6Ƌ~laz�7���;:�Qޟ/ߠL���/V��O򵼩D�lX� è�mI��K�a��"<�J����9�c&R���3���pO�q�a$N��3|�1�h��;�W�<����%� <��"�H�>d�o�;cܭ���a��`Ly6��+(V�6H"m��[ڼN�9�����x����K������4u�@���:�p��Ȣ���@�T�SQ�$��B�y�E�<0�v00A�e��?���j���H���3��æ��`Em[EgV&�qT���YG��*��N�l���1�*��V�e�;�u�h�P��\>��(0Q!�`�dM�(�V`��\1����}S����\�v"#�O�B��?��g�
��0��I}��B�RCOu�sN��dWj�ؗ��
���o0���ę�C,Hd��#����Wo��\]�z�d_��_ T1�R���d���LI���	}�k��L�w�$����(� hP/�@�X�w���HK���лVF��T�\+�7%�Ff�}�X?��}-���8�I�`l���Γy˪%ű/�lG�e[������$Tx��5���a����h��c��K-�w��Q�m�p#Q��W�!��َ��L���)O��,�/��}��wf�?�c�'���F�<����*o ڳ�4�h#�f�K�W�xs��"�]����a���048J֮��O��W���|_�{nW��p��R�W<�2=�ȶ�)>���z�R�'3_I^^/A�gV����ܬsb��,x��9N�t�;�_gkQ^l�� ��}���A����t�)��� 1���i	���/��Ak����\���˲Sy2�ޮ�{%���1s�j���,Y(����&x&�H��m��n,,���;�6n�(N[/M"�;�=�d�w��cJ<V��<I��/i�DLU�C�t����P�S�wE��jQ��#�.3�yܽs�[����Z�ԑ�!(O`�Ȧ�Vj1��w�vJVn���MV�6[�Z��A��P�-�h��{�(��x��ұ��I6��+�W�H8uqg����+�1���C�#�����ԃ�]�$	��6��F$����"e �o�U���e?]M�W"��B/�i.�t�7	4ĸS���O������.%�D=�we�u~7�x<���������z�K(ZDߨ���!փ��d���6y�������Vk���17'b���R���랒�v��hJ�u�]ϑ��(��ȅ�����p���=�*���R����5���F�x�����5kCR.��3�Zn�Z-e��5��0��C���� �okR�����d����P�,�&ͤ��Wҟ�Nz��~�0�ydS:����h�Q���>Ք������g��yk���	�K�kʀ�Sմ�Tb��Ư]�#�R7�U$`�9�]�4S����,��tdul-]��n嚌`�nK�;����Ql���1Xj�K��-؛���s��Z� ��|�������$z��ak�Y��u5�51�U��YRt���%�Y��������K���t�Ѡ}n=���e᠖�&��O� �2�~a�~xg�8�^nigS��?�@����cj�� �iav5���@�K�F��m��b֗`ȫ��'� Z�hڹM�"�,'ȕŃ�Z{YgB��f�k�o�b�m��"E.i��S�4��7�eǬ|[�����ozO�t˛��;� ���Io�Z
;J�|�X!h|Q�/G�/���h��7fS�IF7p�}o�E%�)�C#�=�$M$�|tٻa �ͪ��؝0M/��##����'uAH�4�$0���
>��o0,�U���j��!)o���%k|>��"���ϙ}��9�׮ҷXl����6�$I��S;X�;䚝�ڭ��3�,ܱC�)I�hԽ!���/r�+��(щ|��vi��U��>���n<�[A����f��*&YA�!�B�5��> ��#`(Pˇ�o�U��D/�9�t��JoC�ݬ�����re����LE����P�e*ğ݉�l��(��<�8e�?x* �x7a!R6�!?��f�ڠ?�K3_W��=�Yã�h�LJ�mv�?]��D{��lR�d$:���_FLt�4� *��z�8�<t��"���Q�T�^NX�N5(j����L�[,C��.ԋkjR�8�e׵y� ��\�	 ���,x}>�E�4�����LO>� J�%��В����#Z��;m��-T=��6���:��bʧ���(�{�Z�i����l��U�܈�i�zՂ~է�Ű������A�8eVGI�B�T�{)Y��WF��%���ҭoπp���Ʃ�&S>��n�x[��^\��AW���; � N�?@�h���	Ӏ�[MP���J���gl���5؉iv�!�h	�2�9O���\�Y���1ƣɔ5�aY�D�}@i�e��@������'n�Ԏ�s��K��=�c� [��a?���*�Ĕ_�D�Z�I��Y帮��	i�vv�k�'��;Y.�|t��:�:�b��]�I��H�v*߂[|!׈cw��:8&��e�q|8�tsH�R������|��>ޣ\1�8h��U̍bp}���2*v"iΕ��{b��oWM+n��
wT�:���*�_=�f��<���ہ*�����hwy1�|��u�v�����Q�YF������).X�O������[E?�2�QK�>g�#mu��w�[+��,o���mCf�,'� ���$8��|٫�+@g�H��}�[�<p����F��B8��]�ܴʉ�))e`��0Cs������Iw&�ކ��7��UA�`�ȯ��^��ΎX�	�0C�D��g��HI�b���r	1Z��p�1�8Fz��1��r�i~ �e]�ۏF�ta�(e��V���0	ً�U�
��@�`�2�U��F!�+M�cXNv�w_���A�|��te��U.��x�,mȢ���X9����� �2c�ߙQ��Zێ��m��I2�pv?ֵ
>E�G��Ȓ�_���_�Hq�`�6��TG×u��G�"�LH�q���r�ƐE!����c(�T����&���a�e����ؚ��R�!$�f���[{[r@�@��I.�����DD&��)��닒���YA�k�D���򁏀UxMa�A���M�}�Y8go-K8I�h6�>yb %wC�!d������=z/�X������0�ٶb�����}ftDb�9������P|>��}9�>�aqY@���JNA��0�?aK�4NU�-��k�n�w�1�1���e�[{���L*&c#��dr;�� ��ݘ�(��%G�WpH9�ct�$�u���;�tً,=C-�~�2"pV���'�vNJa��	�cK���=�#���t ˄�T��Q��+�/��2�	�R{��!$V�3E�»��_�.Ki�)w��2��ǫ��$�-���E��4(�10~���q����e(6�{-�
�B��{�,��̨nE~ۺcNs�v���FYؿBXy��h�eb�P"ȶ��1dL���柂�صM��sa�jO�IɢT�27� S��*�j�ʴw\CvQ��9 �c2�`��ڐD?[r㍗3���|��h��{aa�G�S�t@Y�/%s�ӌ�.p1�in����9��*��Gj��Y�D�Z;�+
�|��B�3���4OK�N���.Y��c��I&#@�^�q')3ǌy�����#��D���~�\N"� @��Ie0�vҘ?1�z�{�|�ىm��!�����^h��cJhl>�����hB���)K�F��$Iu��&灖+��Ö9[b5x(�W�r������v���X�W���e�N&:������A�P}�b�yH�,b���}�e�@N2��3�`�`SM7���I�:㛘v �x/���2'�u�3�	{�Ģ�\X�:R�E���l.����1�u��:ؠ�G;�F
�pO��f�:�K���gq���y���l\4h�}��iO��Tx�����"���)p��Wo \n�9=\l�8
�ͼ%���p��x)'��n��X)�z�(��j��$��9i�?ǈȎ�g��[�����j��ug��NU*x��Q+�x�kw�t�e5���{6?VڛjQK�Ka�ݣլ�"�?����� ׷�8�8y�<j�O��食|GZ�ĳ���.�.����	Ґ�Hy��ݔ�Rr���ղ�i�j�V�J5�m���Dr�|Z���c����Hk�":l�ՆI	�p�&0̣�O��x�N����k�t���bS���|�׸E����I��x�[��
�i;q���n�a�OE�s
ݔ��V�!�{�'��4:�7�ݎ�t�0�wa�,��`M��n\�$5G�q5T��I�����'���',��Q�U\��k��I�̆��4����A�>����g�J��.����Hv��|��kㅘyk���षׁ#	�Ӭ��XJ�P%�)�{Yԭ3�5����"���|Mr3��Rk�:��b��ʭ.QrJjQ�y~�%�ӱF��: R��*��L�~Y�.��&��7C(�G!\�;������*�a�{"�?����+9�њ&-)�8#��s�0O�Oaw^�f3�l��ӄ;�v�<����l� b ����3�H���'�";>�����|R�Ltvx9k]V>/H"��mn�.ڗ��9�
��[�������5ڡ���8�y滜#�sZmp�!�{7m���(cS>�њ��Q��(��V!ALS�:�������a_��m�.j�^��m�v�V�o1�l�g�E��E�6#;p^��R��e�V3)�;���h$g� R�CIlQ����?�(7�>�w�ش��_}��/�`C2��&���UcB�5����
?"~��J}y�B�J�O���N m�WE3����[
G�o+0��[�����d�)� �hWJ��\��������Z�1���;dӎ,	Cƶ���U�d)��:|�u`U12�,v{	�F_ɂlk8Ф4G��.Y��bw�!�)���;���V����հ]��p��{&���q$�=����(>	�yr�QrS����Fp��&��W�3���!���/@A8r��d�ӗ����#a� ����	V�s�B��#�#ȜP렫����Z�Ӻ�j�@qǅP^e'=�ۉ&Fv�������ޭ�k���ح�s1��tB�V&��\�#�8�ȑWܮ@���,!�!�s��Z�㢭ž%(����M�ώ�q���'4��|��=�q���U�s����M����1��7�'8Yt���-�.?�Z��ޗ�3�	4�YU��D'�,���y�ޕ������@�t4r=@ٻH@ƒ��Q-v�����Z���FP׼Ӵ�R��Pۚ/=����s]�l�տf��y䍉��R��Z�`b�-
�$�|3��9y�g̨����=�z�n��c�B�I#�vr�1��zk#}�6��mrT�Y�n�BIS˧t.Ten��u�o$S�E��o�뮓Ṳ� \�;iЍ*k0P�鴁A ��.���p������W.e�i���b!g;t�˵CtQED�������I���d'a[lP������C��?�P�2��uMT�r䄈^J~�P���u���K�Aɐ��,�x��2�O�,�5%��M�/�q���D�x,?��ԛ`msl�j�[(�Wo'%2���\}��K!I-��<>��,����oYqk��7c�g�j{��|���.e|d�@Z�_:ֈO�s)#(�{��  �t-ͯ5���^U<���L���X'���
;�+yl��WÍ�AU_r�Mm'L��&7�!/W65�^��.��G�2İ��?<%$�]�&/�24=�P�?�3��0$	�i�ʌ��<?`��)ń����a}˖�O��C	 ��N$@\�	k�Z��m�Q���p������{|��g����q>�V��8E�"�h�S5+����1� �K,��,�&키Xᚦ�J2��+^y�<�Ă�
Z�#�a��������\yJzgЯƳ�\�RR�i���y9�[q��������rK(6�]q6{�2�>���pI�L{6�
��;���ן��-�l�K����|ϜK|���@)B����C�]��9w�x��3��r��I!������P���+e�&NB$o�n	\�]�������)���8��]NN�?3�5`ݝ��-���IR�꛴sl KG��
W"���u�����|���@���W:nQ��S�J�3�l�u"�#:t9�GW�DF�-LO����z��LgC���>,\Pp�}>��O'6TX������t�)�1z���\�5�C��T��Xdl���G(�)C�*n�x�t�?zz����?ö��V���#Ȫ:i�id���q������GUFB�w_<ݔt�du�]M5�l�%���jmq�K��Aݿ򬢾�C���~�*Xͷ��N8X'j��=υi�|���q����ܼ��`� ���:!w	�n!H!ő�i?R5��>i-z!V6�5g�i��o��r����֭[�c�����Fk΁�l~�e���(0�0OT"x��+S=k�/�q���g|��E��І���x�������
1��i�5�� ���ϩE�F
y}��R��=p����c�P�	7n�>�_ރ& ,��M�Ce�+9$��VqQZ���x��ֻ�����,�}`��h��8A��ކ� x�Gx��]��> a˃�$Jc�/�#������t�k�dߘ� ���L��#�����ȇ:X�݃%�����O�@�''a�>��H�r:r��:rn̭Jtyr�Z�m�q~�W"�.nC␹:<$���L�G;�%��3��ư�c��ׁ��$�f&�a$ǲ"����9&1�&I|���\�:�Op�a�����P3��.�y;�%q<�8��;ǐӼ� ���y�TH�i����;Z���9Q���>L��U�<Vڋ�H>~6m
��ڳ*�9�U4�w.��NZC8��=��T��Wl�Opp,;��1���J��iS�'��B����&��MY�Ah�g�֪���+������x���s�zQ�m2U8V�!��E�8�'U�R�����)[���VO7;=~�h@l����d�_�Q8]�[L*(�4l�����x|M}�1Ӿ��A��>��fqfB�����,�
[���Pj}���BH��O�:N�dlWa��nG�
c�OoǕ=u�����d-�.���Wf�#\4 ��M�����1�S��(�dﺝ	�uM�X�� 0��VV�~�1N�-v��b�B��TϠ�þ�dQ�-\v�=�]�~W�1��l��/�qo']���Q����&�{<�d�=3Sܪ��,	2�>r�?�S_�[�bU���^�s]n�P௿��@݁�r�4��o%����1#������Xh��'�Ċv?nP�
J���aZ"�̆qc]^-0=?
&bx燉�ޙӉ��I!�k�pz�ta>sM��t���&��&�E�8�lWx�e����!q�s�VR���������M�ʎ�F,�܏�o���q(�G�q�����M�(U�����u 'T�樻{��Ij?����G���i4�ybUe�')Z(,Q�+yҬq�������fu4��M�WH�Ʈyl��q��'x�q���aF�z�п�RQ�q۶~y�t���)xs^�z��L������5�����`�"�-&�s�Q�^��	��3�`���z�=َNVB�F�#0xǵM��z��R���	�H�uI;
լBe�r���T�����㜋l2��Z��2.���Q��ը ��8i7�!*�a�Y�A��h.��I=���W�� i.�k����;0tU���yC�ȉD{7����]۞�	�4'��cP�I��i�C�����۔���TzP< ��^�5P�vu8���zAe���H6(�@\7k[N��%�i��3��~x�-a��]�	y�����[ĥy���%�r��C��-�II���7�$A��!퍅���/���u�ռ^$�-�����z��=��-�"Z���3���^@CO��p�vۏg����Y`���0KT�<�Z2���S�8tԸjr���UJ�۾��'\C���\���J� W��V�q+_�o��%q�[�wq6�$�*R��^l�a��*��_�:/dD��,Y��(Ss9�޳��8lD�d�]���>Nݘ�����'��9I�,~sX�?�슆	��`K�Ͽ��A�o݅����A�s ����"���<�,�e�ժ$_{�h�.��r z��E��0�E�b{`z�F[�&��s@��OG��l��f�Z�yь3�?n/ψ��d�5�_�v���a�����lX�I^�����Y�J�V�+ݍ�����1ߏBz����p���Y]��JMr�EM�\W��{����ZT��V�b�g�`(�6�q�3~2&M��I�-6�ږo����_�q�3��b�C��r�&iDK:��Lf���H��kADv'/,�X���zـK���_ۯ��mq\��%�8�f���Xc�;}���\I�I`IҲ���m-%������J����w.�<g��
2�g0	���D���I#����b�g�1��v�mLKP��. }�C��;������滔�&�@ع�%=��XА���]h�ڳ�XU�&X]�vs=<�۪Y	{Q�r�\S����;b�����\Q��YQ�ˢ�@&Y�r�z���фox�#�Z���\�ao ���9�ӆl���PQ��U��Z� &�o�ql��^V�"=�S�&�귇���|:���<k���}�sv�at'_�&/�S~�8Tg�WA&����!z�s�LN��D�C߄"a5M����Z~������x6��+�qq}���Qϻ��MI�*v�w��.~Ƅ'}���sڲ@?���\�Ò4�\�UnV�'R��,�b7y;��8�c`�¥��4wu��`����Ӯ�6#��F�����rL&F�7�ӹT�RZ�����cܽ�ꎒYgs��J�1,n�ˆ��~���>���(�+`G4�-��"��)��s�p��V�脧 %�z"���ט`B�I#�x���hz�Ba�;�O�����TSX�B�ٳ��p'T*�����Ɯteu��p*�[����>� ���i� �*�y���*�A�� .��U2��1�WSf�iק�����;׺��0C��!D�ed�e��'���a'��P��|�r�C��&�5C��J��T����^��P���uA�,�˵�A�C����R��2������R<���]�/$�xԪY`��Ȅ�/�[���t��%�^��԰a�v(�I�][�a�<����jѻ�ua�����*g`u� �^�c�2�Ѭ�CJ߹���"c����y�:��^�zC�@�p<��0�ȸ}��Y7���0���ujq����Ng|���S�r����J嬋��w�1�I�Y��8�Jթ;W�
wV�:�_1�k�?U�Ut`w�[g$�ï
�l�f�3�?_�=cd�Rñ������9+N�tp	l-�b����Z��Ꭴ�X�'T�9�~<ve(dڊ�����
!�e�\eF��m�iS?�
�� �\h�+N|��1�b?[eR�$�h)�c�,.�l� c|"E�ej�nE}�ǛzH��[:�O�Gp��q���j�o}:ǢQ`H��rz������I��KI+B��������4��L��,��ԔXrF���:$b�����K^y�' f=@�EP�.����$�����d�s�i�+�{�2|wS�.�9��@��_US�<�t)��{�U~ �lA�'5��OU��!��bg��8�6�^h�y����;!GÚ�3U���.F'9(�&��/����O��ĵG�f��~�D/�<>�]<]�/�{l4
U�E���^	6����<,��Y���V�.i��?�����	�s�NqJ����^Z8r��~��=,5�+{��èb�yi�C�n��FO�O�chO9�5��[��B���j��0��Ѻ�r����c�g	UJ�\�+kM`��q��$<�����mp��DTk<�J�@��Ӻ�\�;����Ӥ�A���j�m�pm��A�(CR�q���24:���\IKO�6_D}F�Z��_���qb�����RC��q´I$K���Lt� ��F��y��//:��X����hGKA�_�mET���\]|%D�f�u�X1��}_E'��In��r5���@�%7�#�ѕ�W��ZO����YH4�����{���!c�1���-H��ÿ�GEQ�䭐SI�� ����6��M�O����ز};��f��ǕH�g��f|㫅/*�����)��gf��K��x�.��z���Da��쳢߱8�0��vr�%'7�2��-�@� ����PR�u0����K,�[���R�V_��^akTg����������,��?��կt�����J�g��l��o���3��A���9�stry�Z��`�i��ῦ/��Aݯ���D�?���i�a1��m�j�*[�����ޖ�(���!�t0X���Vm�A�,^Kn�^�6 ��(@!:MH�v������i?�c|�d�!0!�c�?�6���u?j�iT�P�>��i�.眰����3��ܯm_���U�f	1�C�J!"c`�9=����j��iZ��Fn��M��6M������֣�{Ե���D�DJ���6����H��*gY�����1�੃�ri&8���+�]�7��Q6���+��s�"�؁!�Pꌰ?�>]�w-"���/Έ4.�v;7{|���h��t��Od�������D/G�e���7`@g<j�G���$s������eD��3��G���m5�Y�(JO��@�V'��#1jb*&�������|��jѰ����C%����O���V�fF\pGp�=��Q�f��9P>U���R�ԡ�p����kR ?�3�e���@�hoX�Ղ,��2��_ s2JR�����R3d�c��T�����j��X֤ ϙ�pՙ0�WJy�|k:�t㬨|}Q�n%>Gm���<tc�g�.�y݀����^K�QʲbSG�fT%K�>��r;��o7���`��4���S�KwؕY��rBd��-�W�n���`��d�mi��y�OQA��#�;�}L�-JS����Lr6�R�z�����;��$�VS�u�|k���~�x5#�����3YDKn�5���#�4������u��.�^����n/���,��D�&r#ٳ��2ώ�������ɲn[~7Ș���ڟhQ�ȷ�%i���"a@T�}83�̟n���h��I�qȝ`��Y��Z�"~��U�"�4�^$ȕ7'�Z-k�g4�hf'��oO��$�"7Ƈc�4K��k�|M���o쭙t}������ ��I�FG
�8|��s!���:���?�Z^7���I����D����[N�#
@u$1�%�n��L���?�s�2\0?�����#jب�
�u3�e4|��I#�>l��0��U�����i�!�y��z�Tk�����9�7Tϋ���k�f� �X����r�VĻ��u�;
��䌣trץ*k�c��);��hKr�ґr�p��� ���wFvۓ�U���>���������������LXA]���ی�AV>��I#=�P=_ioM�6�D9�n⋌�[!��ݞ�$��d:e/']��i
�� �����*62��aM5����nvaeb��*��+7SAb6 @ ?bj�����=��W��F'��l�L<�im���?�pD�i�^�_Ж�����)*Lf�2l�����
x��O�ISƮ^���@�Cj�3�&j�U���m͋��s�����g�t �>�@o��m�)x/�[EzE�)�?̈́� <�e%�=����Wp\Z���;�0�͟�����~��F�D�T���(kZ�Z���Y�lk��?�2�[raմ��h�Ƭ�R�����8�����TIB�H|�m�0Y'dDFn�%���}+�o���HoW�[�=S0��ҠA�[��\�w{I��m�� ���?�hub	S�[�*A��^��� l�H�5J�5vsQ�h���k3��8��Y��w�� >�?v5M� ���2a��[�5���� ���$'�̮� �Ns�;���=1luriN��a��X����6�S��o������{�_��zvh���Y�2�a�.n􂻏��:��ϒ:ĪI�v�i[�������ABм�`q9�}Àx`H��g��*�	���+��U���*z���b��(��$�*hݳP�7�jH`b��aoI1^n�.�w�0��w��*��D����<u��3� ��V����w�+�|]C�h�i��Q$=��>��̇)`�|����I�.�Ì�?"�vQ�=r��J�#_�����q+�y,!k��_F��^o���W��8t�2��D�+�W����}�0�<��%��F��58��]�����a)���{�hs�#��<�����V_��W���T�B�x�Y�i���V�d�5Qդ����ґBOU֗��c�M�� �/kx
lh�K���v��0�� O>��xCsa�8�kQ����i��N|���Ed�����x���p�
ۗYi�g�*�%�g$�Ew(�
c�� G��������P$�z��7���:K����0,�M�4�m$��!q{��Oa�������>,��[�.�1�ȝ�-]����*���>
V˭=<J��9ӱ�H��:n��ak�z�?*���F���?��)���rV�XЁi%7�_��ѭ�������h)l���r�J���{%:.�����&r�-���~���P;�ȭ:fY��0��L�oX�8ܔH`9�=�m�R����N����[a���"}o�:�J9���&�r#���O�W+a=����n�3�r'�颋;[&�<�N��e�8�&DD ]�c�fH��-_s;�
���Z���sLz�g��=V��Hh`�mt��]?�9�뢡B��&��t]�'n�~YX��]��9<�pZ K�����W'�u}�S� ^�9�����VO&�7��A����@lɋ�Ê�'?��O�4w;�$�pm��V妨�r����e�?R�|�hv�tfȤ��VyF�;�rh��p�����jQ�'ƣ��(�P����q��:}t�������\���T_BG����
�q�ٚ}?q!B2�GO��NWy��X��
�Y�o1���`����dW���&��W[�\��E��`�\1�3����dw�	I��������s=���{d1�j�v'��-��r���G���Ͼ������e�GW��f�����w{(�[G0])Y��R`�Y�@&y8c���=�򥪠l*	��r؞~S��Z�'᪬e���A���I/�L��@���r�u��3�p��#�W.�{���8ǿ9���t,i�6P�∙Vg{Z��̰2q�Zk^�ڜ=)
�&�uE����}y��3�k���(�s�jt�&�&�v���#8U`Wb�؀���!�BsX��iz���wM��J�{���&p��Cmj��qg�ڛoq����MJ6��\*�<ߤ4'�f������s�T?����_���&4&$U��'�66,;n�y�[i��
d�6�ƽ4��|���X`9��?ێa���Ms15Fּ���}R���`oo�^�e�S;Hs�H�2���T�`���Ւ۩ `�r1-P�%컔Z�tR�������2����z���x�B�#�4��>�z�z��|�#�s��X(��;B�Nާz}�T+Sv������R^�K1��F}�q���� b�i�0*��;�/��A&L.J�B����y�W4|i�2*���h;ZnL�PC:�'De�.�&�9��e���'�JJP�i���Ck�T����	�T�����^Г!P��u��h�L�>AO���rIዪ���`��wE����x�͓��8s�P�0P.[�*n��	   M   Ĵ���	��Z[V)	�-��8�d�@}"�ײK*<ac�ʄ��I�`� Px"�f������̌�M�7H��B	w�4xl�9�M�սi�
���L��C��o8�Bœ�,�-���ɍef��A�iM�R@�O��1�U�X<jq�i/Ov1�bJ_�b��U� !�Q:̎�c�F�>�ڈ�t��}�Ĺ�r�	����	'�MK!�j?�?�7�@�^�T�%i�l0�ٚ�
�kR�؍u�Z1�B�Q�ɧS��!���9|�O�B�Ú�|�D���><��J���Ij��n�����|BHB:��l�ѥFL!v\h�m1�yr�Y�'��$Fx"l�(|,(�ZF
��4f$U���*�n#<�Re,;QT�9Ĥ�p�� ,��E�T@@���O�8s��䔑��'��|X���cV��HK�+J��2�4p��#<q�"�3�>P�&%9Z�m9��V�s�,���f�[<#<at�>?�����@�Jqc�hޓ/�XU3])���&s�h1���f�9�*���UIKM��툏���4�O��a��<�м�Ro�,w���"JӢT��<��,�%{�O���P2-�P;K��4��A�"�OlX���d����5�^��	J�0ձE��TN)�m��h���#'�����7�n�� Z*O��0þ��I� @�y���"'�$P�,A�L���{x���`f�	���	�a!��Za�P�RBφOt"]�������׍�5Q�Q����I ff֝�S *l�xĨ"==B�I�T��  ��� 	��v���b��n��2O���/�PHǶ=W[
L|7wCof�p�M��IU=�I���(�@s3��E�co3u�[�7������LL�R����sW��y˙Fe�h����IuHU˳� �{Eôe0��`H�w����(Je��x������:�=����*g$�˭���g��Nj�"�,�>�k#\x���"	�ȵP]E{�U�n���7����Svu�]�R�(H��+�E�5�Xg����#��J(����@����d:<�f�x��IS���MY6��!�
��a&:�Lƿ�1֋������i`��:�6s�K�X|��D�֬ZkH�(҆��7�E���?��J%���J?w��H-3�rL��U(K'l#[��S���RW��d+h5FI�&F<�����^�Ս��z�   >    :IZ@-�nkZ��&C�'ll\�0Oz+��AI��e���X�'iD��  ��K�c�x���,�]d�G�6=�   N   Ĵ���	��Z[V	=��8�d�@}"�ײK*<ac�ʄ��Iڧ`�\xrlgӤ����O�8�p�L�r�D�bBD�.8\��nZ�M��i�B���W&Եz�Bָ~ܜ��I��~�b��	Q�� ҵi�*�����+�d1Ptg�[���+O���a.؝DJl!�^��kI\�bN)хͲ>qǪ�n�KóUp^ݡ'/ӿ0,�$�N�l\|6-ϭ;��ē�[�p[ڴc��`�O]p�plˉF
y���ۍdZ(䁰�݈��%�D�Raљ N��$���a��
;3p6��ӹ��2���~)Ij���;NݤL�2�|r�D�'��-%�\���[�:LT�CHZ�xĀ=��c�h�C�	M��� ᥗ}T����GĽSl�1s��V*�O�ܲ��$
��ƥC5�EځM��f���Ƈ�a��"��"<)UD&�ɬX�|�x��܍L����Q$)��7-�/�O��	����CA4X�%/�$V�Tq����t�r�����!�OZX��OɆ
�-)�T�s�> jJ�x�]��P!�I���O~�����iv�B$�U$EZ(�c@T4Fx�Hu�'�r���5�DD���fS�HX5�T*A+Jb��[��ɩvT�'�<B���SӺ����Gw�D:�'��aExRn�O�	(6�����RS�U�ԡ�]7���r"�*u��eU�h���).���މR�"��'I@��"�5���H�DC�K$%�屧LȹZ����-F�;�剆C��),����B�X�����ٯW���2Ѳ]�ԭFy�@U�'�부'�$IAo�%([�y��'��@ ��FJ	l�V	�R��^R�# �A$f�$�$�O��d�Oʓ�?I�}�d�3zH�l��I�W4΍	����=�|�Z��"Hy♕Vn��� K����'������Dݷ*'|y����	K�]�������
q,��P`�v[1OF�˦�#}�oM�W���&?!�B��q��%�+׆H��Q��*,O�R�`�����`U����p�Z���7O����	���D�Or�2^�� �\��"��b�1I�}���?������O��fD�A/�arU΋�_��ӌ"4�S�4M���1��M�F�`�I
w���x�'�qO���P/�r�'#���Ӗ7<DZ��ҿb>�9�����<A2�;�V�>�O�Q"���Pc��C��[�$����"O��y�G�t��5���2D��ۢ�$,�S�'_\8( ��$��Jg�/I�8   >    :IZ@-�nkZ��&C�'ll\�0Oz+��AI��e���X�'iD��  �������T <�<�o   P   Ĵ���	��Z3Tiʕ.��8�d�@}"�ײK*<ac�ʄ��Iڧ`�\x�	g�l����5B@��"!HkP�����L�TP�PnZ�M��i�����Z�:r��
��9~t�ش�K1p\�	���	
!���Bѻi����	� �0�ҡ�ȏ-����)OJ8��$�*#>�x�CZ���
I�:�����Ȯ>`a^5ehTv����D
ӆ2��=��囹��N������a����S!��)��~�q��. d�yu��̲D�%�S��P�����S9y��<ݤА�/Ƨ	u���%u�&Hp�� %���+��U8��O�Ӊ�d�����e���
�v��N#n����'V�#<��$5Q�ȍA )U�j���S�[�t��)��0��,r�Y��PT���u�e���ǟ^�|���0}��Sp�'�P��=Q�H��i�x�j�G@�*�������5���	���Ԡ#�P�-�K�B��0��hVL
8e�Bc������	�k]@�9#�E01��=(��;5˓i�:#<�1�'��'`��@c�Eԙ�X��R�̿\�̄��I�0?�����'"E����XϺA��$,6`� �yb[�'7�%���(�H%\��%�)|jY�Â���)��7ډ'�����2�bX(b�_
� )�"H�P�V�m2w�<	��.�B���Mb�õY�h!�'�6�;z0)E�� �Y����nM�'�%��m
j�''�\�O�8�0鋣=�,��p�;i]b1��N�./~0(��ɼB����DD�M�� ��'��I/��`��9D�(��*   �z��yg!>Cy�B�I V�����ΘR�
 б�0l���d�U}��?ғ��'��1�1,V�y�hXs�O�]f���'^�6m�>JqO�����^̧7K��r�Q��8�*�q�xT�ȓ
�ɨ�E I ��TB�!:0�L���y㤘�F�р9�(�'��-�Ą\�}��`��Źj~ʀ�ߓ+��'Ir}@���0os���� ��䩒��:��Tig�'F�Y ��>qh��'�j���N�X���_Z�b�,�e$"�)��\W��9(,X����N��s�!�DG�'��a�3�j�@h(Q�Т�az�$���!s����^�I��=�!�ͳ��x8������
T+�K��O��Dzʟ(D������<� p�O7�H��WK�'G8���)��'My�i�+=�|��͊�o^��q&O	)   >    :IZ@-�nkZ��&C�'ll\�0Oz+��AI��e���X�'iD��  ��ڈyR�)�ӈ�4�B�U   P   Ĵ���	��Z3d)�;Q��8�d�@}"�ײK*<ac�ʄ��Iڧ`�\x�	g�^�mZ�Z�xI�`eS�z��P�ٚ;>R��ݴ	�Ư��!���ˤ�z ]��̝>���k>^Ҁ"<�׫eӬ��re��m�4� ����7�=���R�`�����/ފx�剤�.̣�,�};���TP����p;g�y&ތ�4�O�u^|�m�bG�h͓%�D$��k�@p��?5�!$�+!��ȃ�0��,7�:d'��j�'H?h��,�X�I�*Z�*5�	 �
-���4=Q�NR�J������0�0�5�c��'T0`Fx��y�I	{Kp�iZ�h�F�S ��4gD� e����	�c#��as�ڥ`0	��+�1�&����D�$�O:ia�O^�Y���X����V�Vx��@�>Q��8�^���|�D��	nZ�rG�V�+'��;��y�����͢�O������.�6�X�(Q7bmsS�E�;��O"����D$����X'�b�K�
�hc.8��Ia_�����$�3e$O�Y�t����&r��@�������O60��P�y:'�́�� ��jД#7H��<AĊ/��O�@�m�R����L1"S^h���O������>�ē�M���;��<�Dfڍ]f�Q�G��%�n�l�(�Mc�'��6M�O=�"�����'�ט)���U�U�.ء��&Ml�9�'�6��R��m�'jN �O|�s���lC��`�Ǘ5�(1�͗ ��A2Q��Z�|����$�~�G$�Y�����>D���qi   �k��a�m��^3<d��F�!2�-�&�ο'a��Ex��'�<��7(��8��T���?i8Œ�'y<P⒡
jE�6��22�s��N��ɇ�HO��&��s�Z�R�Pthf��E���*&��h���b��5�ɔ	,Ȩ N(�D
02�(���Y��Y��_/,�!�$kx�9�$�m�&����g*!�dD�e#tPj��K�����@κux�C��f�r�U���!���1��j���D�d�I�Q_� �� -�*$��'�
i�Z�@���D�f���	$S��C�+��U"n�$%R��'WX�o�v|1O�Q���D�^�u�a �늢z���(3�)�yR��)��!�η;���H�)�-�0=�2CO�R� ���	-0�	���y2��G�N�2b
Ĭ{�0�uȈ6��'E�"=�OLR��f���eZ�   >    :IZ@-�nkZ��&C�'ll\�0Oz+��AI��e���X�'iD��  ����|
�  8El*2�   t	  �  �  �!  �*   �pA���d���\�'ll\�0BLz+�\�u���e�2b�����/\��'�� ��f@�T����B��Lʀ�Th F�!C�'S��ȥ�L B���dC�lp�j�jƈ)��'���T$q[��Z!�557r��T�J��?�����?I���'it�I@ =��
��A���D�	�!�'Y�1�0Ɯ6����E�s�R�r�{���@�r�+Ib��Ӯ3��a`�s�@��5)�\�'Z ���$��'
���J~�3��k ���e�/m���Vk�N�<)d��aԀ"�FFuf����@�u��@�?q0��/R��H�Dջp:�d���\�<9�T>;�LL�b��2��|����U�I����hq8���t��������i�鉪c�$8�y��	��zQ�t�q����D"�"!A���'��5��k�g��h|D��D	���%{�+��rC䉘6�.�[Sd;���Kʐyjc� D{��t�8�<X��U8tppьަ�yr��΄�34�C4;�!��[�Y���(�O`�� ʄ�	o�� ��B�7~R��� �OvP�B�o̓yQ@F�t�ǘ
i,�br��t�N`�Oµl�����1��?!&�M>2�Zt)�����sR��r�<�I���,bpOtE"Q�q�'e�yR��j2��!A�. �&��˄��y2�84�F+�V�&ž���"C��?�P�@0���	Y�I�[V&]8D@��r�t
fG(��E+�e#��l�B��J���2�O�OT��©3�b�)a&V�b���u`��x�|�� ?t�Q��%)��hE&A��ļ�D��>����-,KFF��-����z�,�f��O`�d�Od��<����'��d�4���Jt�aX�-�$��3"�';�r����&(<Zb�T�9���{�D i��P��00�1f�O��Y[l�:6��l0��)��tM��!��E�9��'�2��E�^y�:)j�A��ݡ38>1���G�����d�&r���K>��OD��^�G�6�d� 7�XX��0���O�$�>I��ɒL�M���<��(k�P?���?���t��:2��V�H�������ڦ��'E,#=�O��eA�l&+�Û9�	�S�T/�\�	Iy����YX�k�I\�|@/�;6�D�!d��n�|��a��o��i���#1�ɫ~�q� OF�����L�Qg&I7KJJcS�x�+�
�O�����Se�(p���"&�4�leSW�x2̀�?����'�ħD�`�	��6qY$�_ip*`�=����<A���Zl�	�[;o��N��HO��Ӥ  �㟼�R��(U���"b6�ֈ�B�(�����?Q�v�z��V��?���?��<�$�He�΍{#�I��M��w� �R5m@�o4�p�O��Y���#��|���fܘ)��аn��BsnF v#�\�
5}���y�b?O ��� ȀY��Hb�O�E��d�ӟ���ɟR��	��>��M����Rm|�v� j�4�g��
!�䓰4R��)$bF�@�Y�ր�!b�r�`�����!�uG��O��},PЪ�..A��$!�$�8>��`ڷ�L�ʹ�'��T�$�;י>	��\�Fv��e�� ��wM�O���()`�3 ��B��Dy��������;D��c̩lO&�9�ݰ0�Jt�6 ������w��!�W�ٻS)n��b�ќu+�ч��.ܜ��O��R, ,����F�=qk�?��B�h�l��	�"�iӎ�J�(G/*F��ǒ'�"�
6-�OR�$��?4�qĆ�O��_$tj&n��I�,@^��vɝ�`)P���+��V�r�򄚠=��O�I1��w�v���A�c����0�'������?I���M;�e##�v ������|�D��S\�ǟ,�?�� ��6���:�jD�~���2r�Z�r^���v�h��WA[&�`낏�?w�Fi�.ʝ�?9)O��fJ�:kU���O$�')o1�ߴbD`�0F�v�HЅP<X���'r��7P��c����y2�'��t�a~re�#s�l��D.��sJQ�䯄���!D(��ΛJ��,ݣ�h���a�D[4�A�R��R^��@��x�7�?9��M��'Ա��b�ߨ*�����Y�E�%�$�O �=	�O"Tr�)ʏDlػ���	��`
rE.�����>��x�N$I+�]
U�R�k�aq���E�@��O���O���o���D�O<�D�O��!
� *4c���	Ue�2 ҭVA����DȨ]���c�=�?�'�#:#�0��&�L<9�.Ĳ;��e�Ro�&Cz�90���#����1�����M�:�p��~&�D��j�-~����B�	u	E��?!�O�0���d�'n�O�hpq��V4}��K�p�qRV"O�u�è�dQ�<2�F�{AN�"C�'z��	�l�\#<yTc��<��OdQ��Gν`��1;�ϔ�|N>)��B/iA(x��AR���	՟��	'n9P%�w	Ο�̧H-���N�s��!R��A:_*��Р�a<�Ĥ�5��@c�-M��t�����B��x��4j4p4=�\(3���]_��P�ӟx������Ixyʟ�'�B�"D�C(���Z�/{~��ߓ*$�'�l�SӇB*s�}b����ɋ{�`�>rIRS��RB��!P�Iݦ��'�U[ڽ"1Y�R�q�#mQ��d8�jK�6R4���l����2����<a7¯Fq�$qPg�3c�n-��d�kX��@�F�=^�E[s��c����"��x�U!�,Wn�9 װ<� �����	��Ms�4N�~<�1Hׂ$�X�@F�w�~��4_���ID��|H<1SB�2���@`I��rL�M�RE��.����'m���%-�9j�KY3|�t� �o���?)�{�lʥ��$���ں�e�CO��L��.Ē	_���p/��ޘ'�؁2uO�V�g�tW���`�ρkΔ����'��B�	�>PP1�e�\p^��NU]��b�F{��t� R�6�5�]?wX��+�2�y���X�$���bX���M?B:��L�OT� A�^�e�|4 �׽r����G�OT���!�|�GŰ=D��;l\�Q��nl���)�$)�l����?��mO�eSt�U. &�-Z,�v�<�HƁA������<sf`�S�KW�'�y� �qj@�G)�#o�v�Hâ��yR,�;@ynٰ�F^�;��%��f��?��S������Z�v����˅B�dT�r`ZR݈�	!0���I�L-�	�!��q�/!��L�X��	Pf�]$W�P�%��m^!�6] \���� :����Ոt!�D�	!i�U��`P��-eǺ�-!4���%BU��4`�V"�`K�E9|O��'���0�ҽ5�z��&%!:à`qC;��!�HOd������C�K	��1Bq� bc�ȓ�4}�җĒ�3�y¦���'G�5�p�Y�f�|��C�&���v$L1��V	#����ԯ ɂ����o��XQhu�2�0q�90sM�|9�D�ȓg��LzD�X�I�DԳ2Ć�>��?0�)*!EҸGD�hc��8$@�K�D�~4��0�ֆ1ܘ'Š���'�FQz�AI�\ ��`���:5Q �a�y�`%"Q޵�}&�x�,W�%#�A'S����>D��Ӑ�-"x1�)J�yݐ1���6�o���O'�4�b�P�%{���N�\��]��'�PR&W!��9EςXjPq�Q�e�ԉ&�I���A인Gd`�TO�4�T�Dޝ`; t�<yG�U�O�eI2k�@�x��Jl�A��d�r����5fŻх� 5!L���iՉ(�����2N9I���!B��m�$(ޅ&�B�Gx��'�VT�C�U�_�P����1��'2,�pR�Ȝ2%"��`�7|:H ��[��ɝ�HO(A&���UB��ذ@�rlL6b]����Ĩ�Pp���+�Lb���Iګn��O~*�H��7L\1vC�A\���1"OBm�a��<�6x��D�=K!Q��"O�ʓE�6���q�*Z�0<�u0S�,4��	W&�+�(��"��V\0ܒĪ(|OF�&�!e�7������i�pI�f(�	��HO�x��W�2��lg�BA�4j��-��G&}"����(�y�&��'g��-v䗃-��q ��(-���qK�AkT	ϳM7 P���/;*E���[��
D9���Q	^2ry�6����ȓa}�z H O �i�B�� 2��8�?a��)�靉z�e��٭ט$��W�,d��lr!����'h�uK�'mּ BT�ĘaB
�`����z<��y���,�
��}&�� $T�a Z�c(�u�oP1"�"Ox��2��UdT�'ڢgif0�&�)�S�'�sR�
ݬmY����WЅȓH�d�h�HN|��٫d��8�R��D�|b���жL�E����6����ڹ��ih��!�2��Rg&#|�C�W1����FY���	Z�-!�xb �BQ��Tæ�0�pRE�Z�[J���a&D��Q1�W�k�f	�g)^>aL��e!/���<��!��YX�pǫ�8|L��m�N�<!$`S#3����1�³��c���ǟ@X�O�Gz�>�$���;a�'�Rli�mʋ2|�d�?]���c���[���Q�|r�ڦo����5e��|��5�Eȃ��y����?�8��R#�h�&�
5���y��7A^t@��+�0Dq4l]����4R�`��9SP��!��+h�{�@:�$� 1����0@B!R+Ќ]	�O�Gz"�3"�����4K
E$� ~�L�gC�4��<T�4*䣂a�4��A'?��ńlF �âq�%��"D�(� ��	=���/� *��*LO⟔q�/%O?��h� PU,
p[��(D�(QE����),4\ ��� ײ�����?�2Ay4�zr��-r��D-��HOjIb�lYC̓�(!�S/3�H�-�D/����N�#h�XD�<��B4h���>�O�|h�#ǊeaP��M]�]�9�"O���S�K�0Gl�)����0�S�'=6i�5cM�sy�]y�� ��l��#�$�Yw���tÀ�9��^)����|���/[,�m���/I�2��m�N��f Bb�4k%$%§М5�AhT8� �M�b=�hs�O��P�`Ն��a8вo�8D��pu�)\��C䉺zԌ��ᆸv�جXЬ� sC�#<��/ה�s��Ҹ�J,(dN�3�����IyZT�bZͬ���XK*��	!��DAj�'!OΨ��#Q$&eNjcd���X$�OT��䏤\�1O���!�Okb�'Xx�K2d	Y���d��!Z�J���'��� �יT��1"Ĥ�bհ�'����ce�'j������0K��RO��)�)+���Ff�gX�X��'h��Od����R!M\]#��	#mƊ����DO�'�zD��O�$	P	{�<�pa��?4,�U �>��'#"�<���l������ i������7xU�B䉦WV\e��ƀ�RM���5����<��A�����W�:5ꧏ[�m��C�I�s������ƒw� ��GJ��{׺㟜y���?�X`L�??:0�V##
J@c�l�.�HO��ѢP`�8Պx��`�|}�"�M|�����M��A�<�WCLM/"�>�O�pCe�	6>-���e�6$EJ�a"OX��E�˄^�(��F�Z8��P�!�Ş<m���K� #ߺ��cG?tz�u��\n���F��ɊHyGM�=��;��|�f�DD�"���#֣:D<�J�Y�?Y�ȅ�c�,+B,<§�=����'p�-xF���"�,��i�ԥ��I��.�v�7 �@l@�8�LB��!ۨ�:�I�9�8��3�>�"<�
ϓ;`z���Y�2G���cֱT]�Ї�KE$a�Ф G6��� �V$@��5�I��DJn�'��OR�B��Y�hF�V�@刀���O�I� ���mI1O"�īD<.2�'j@�F�)6���*V�<3��԰�'�6Y2$�E]�R��%+8.s����'��+�,�'}�Ĭ(�gM,����O8������,n�T�2i�-�2d*1�'SؓO.]�A��2�ׇ��)��l�$��}�'���	��Ot�b@�</~J�	� J�q���>�f/�\e^��<���O�3<�-ha�J�xM���!3Q��B�)� ��,[�4:쁣Kּ.R�Y�@�'�O>����HI�=�vj��ޜѵ"Ox��a�h�Āi�I�8��=;&��N���Iǿi���6gέS:���`�Fz��c�L�7@�2��ȃ=@�*�	Ԡ�|�*7�%扑���zC��|ₓ6���h$*�q̣���<�yB _;99�dӒF�5ߘٸ������'ўb>Q)�E�(Z����4/���Z��*D����E�"p0e#���*5��5�K�';�S��'j�UpkƣP� !C�(�V!;� ���2��8=>=VG�
K���[MD~�&�!�IN3��H3�?�O��z�KJ�j�G���^�4�I�"O�� 0H�	S�X�X�Hef����Wx�ЁW#1nH�D���gаPCw'<D�L`���g���b���9r�$��O�`�'u�"=��|��S3h�y��U�@;�;0���~�!R�!�y��E#R�!H>�#��H@�-Y�)K42Qz��d�g�<�oO{��i�s%�<�Q:�C�M�<��e](czT���@?�|�-���x�F�.3?
с`o_�pTFժ�E ��=I�|rL�;�m"%�?f�֍j�	"��'��#=1�h֝p8"��5v�� �I�n�r�"4�A����y����G�%�I�����>�"A G� m�ڳ�/N#�("Od|�v���ܛVl��j}Qf�'t�Of����L#�9�P��eZE{""O�)��=r�4q3S�VHx�"���B���i�w��pb���'?2�k�+º!f�ɖD���y�������G��=��*���'d�-R��Q���'{�tᄬUm�g�	 A\(����ٝU�,q�J
�D�B�$Ig>I��'��v�B���F�?G
b��F{���� �ҔR�H�F��Pr���	�y��0tl\�*�ȩ7v�9�f�[��ؗO>��t����#yv��7I�yN,���K�O� h�(�a̓dw^E��[��:����5V�Q)�L��Otd9B�[��?�@.�1<®hBFӷ���4F�<�6_�1m���)�(e�p5B`L~�'��y2��2��Iu� Q8QqB���yBD9;�r�!��-FT��ֆ�?I�Z�t���p�	�dl���$��iys��/z`�	7���ç4所&��[%�&�d��OP�P`�+PqL{$Ņ�L�!���%�N��֮�<86l�$�o�!�D�&(��}���]6��˴#��0�vC�	#g ����(vg���$��$�����q��. mN��/�݂��d!��+0*�(S��FT���I�'>X@��aD;��\���)�
�'�(�b֩���'�R\�O~�qB��JA7��}��%��4{!�� FL�%UDL^�!%�ƣG azR��T	�!EF|�	�F�<a�!�Q4�h��N� jf�IB[�UR�On�EzʟXa���=�B��b�t�쌻e�Ba�'�,��?�I�G�(�I�g� ���ɓHs2v��IQ�`$�	5k�H���|���y�0p�C�!4�\AS����y��&^BQ� �&"G�lQ��X���'tўb>Ic�"�>�5�5�
?;���"7D����4L���H���5�)h�͟[�'�����'w��2�
&n;R)!M��^��(�<�^�A��IV>ݘ1j�/|x���Y�R�sA�M" ��96	&�O�i�����]�	ւ?p�b�"O |��BI�^
R%�E�'���R�	Yx��@�'��Q�J��qup⠈:D�0{&�N;%d:q���\ _~��H�O���'�J"=1��|R�y�0u�种=� ��#��~�n�7>�4�y2�L��F2L>A�C�R�t�+�-��14]9�Z�<!�_XĈ$��.��QS�X�<� F�K1�z�Đ��B0l�p8D�!4���$A�2�@��/$���D�%|O��&� ��=&������.
��K��7�	:�HOXp�Ul����sF�ߑ;ZB���m��8��4}A�f�Jl��y�I$��H[X���F�H;�� 5owJ8��c�2���(ԉe�
��䊨PȤ��b�q��B�'���	�
���ȓ��Qh�o��t���[I]-�H8�?���)��noGZ����6z<0���a� Cߑ���ǎܘ'ql���'izz��	%7w��SƝ��ʏy��	/����}&�h�@h��?��`D�_�v��)1D����	��{Ѐ��<Eo�a�F-��O���Oܪݙ�G��斌]`���Clߍ�yr"W��AjNT�b��kE����(�O���[BJ�3
�ڡ&��q�Ax���%e����T�?��Ux�N�!���i�O�D�O�-��xa�aA2}��I�A�;G��L��!ܠ��+S���
7+�莉��~&�`ЗI��n<%ץ�R�L逃D�J��I�UG�F:�(��'(c?O��M7v���`4���tͳe������' �5���|���[�C��9V��Z����=�!�S���\��*�*jY�03����!�mc�TY��?��?j�����?��LbA�S�Hy����P~h��"H f���c+�	K$|��3#}��=+w� �SE6�����-1~��� �S�xwEħkV�y����IP�U�9<8�s�J�s��͛ ��3ņ���eϛ�pX��	82���B��8�F��G�o���h"�On�D2ړ��':&\�T�6i��xl?b$j��	ߓ|��'�p� AX,���)�M����<#�{R-�SD2W���'
5|j�Φ�k�a�e�E��MܔM�*�3�, ��?��Bͮ�Q4�1�?��OH�I-=r�j�v�2<:��6�
��K�#2d�@��q8��J��7n��b��&	�q��v�ḻd��M����4�ڮ�xB���<������=J(`�@B�H���PRm�5�qOt��$[H�hIu�P+s��ѐ�"��#��O�0Fz��%���4_R�����]�貀	��� `/J�d�<��M�R~���"H��?i-�*��g�v�9����	��8����h5 PH���1�?��a�0��FiǺ#��;�FC����_��,Ca/��?��9b�TQ�!�$�L8"�9���Q�Ș��F;$�ԍx�J9�'g�T9; E��r�����ǒC�|%�k�a�O��$>�'�M;�M����EHD�\�/dm���I�<y,߻dy:D�uHO�8��d�eFB+�HO��!qrp�GJ�6Gj��1sꝱ)�~m*pEK0��e�S�!�?���F��Y��J��r���?��'n�I��V� my�k�*�H�r@Ԣ#�00B���`�Bo�<h��BA&Q��xiF;[qb���n�����[��,���ʑ67����+N�=���L<Y&��e��m�W�Z:Q
֭��"��e�b���Cg �O��:ғ&�Q
i�1��4_���b�Q�<ac�*r�]J��G�>��� �ǟ���'�������O�~��>C(�))H��!�	1C8A#�0k:l�Q�É_�2�'���'-�͠7n�A>���!KEv��P釄�z�$4mQ)*ۊ`֮X)�l��I4���B�&�y�Pϊ]�*��C�;(
�a�i���=Y7卯p�J1���A����⤪�bn�d��ϟdD{���S=bפ��1֊Q���seO_H��{�<��Q�Grh;��O��DY�
�b�qOҬ:�"�O���irE�����cǶ7�3�� x;"��.�u�d��#;vĲ���:QI�OɂH��	D*y�p�1(R��'ǒ�C�%�T ,��R�0��TH���'�n�頋[�OK
�YCğ"$0�!��'���S��T�q�_H��V�%��'��#=�O�r(%n�+���h0L�:���á�+ғ&ljx�@�D�� ���9	$郒$K$K��<`�k����'<�C5�\U�d���?IXDAQ$����G)T� �w'�I6|���AX0�qئ��9�S�'`���0��>X�3�b�M ��4�~q����7R��E�(3l�P��D�|���$�(:��&� �h$����~���%�Oֽ(E@  ��   �  �  �     .  �;  #I  �V  �c  �o  m{  ��  ҋ  V�  ��  ��  -�  o�  ��  �  ��  �  w�  ��  �  ��  ��  %�  g�  ��  }�   q ;  H$ �, T4 ; OA �G �M N  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}���'��k�n�����(0�ɻ&	��D��+��iC!�}Ж��fj��$ND�ȓ�v�,�.<Pl�C�k�7$�U��k_����c$�I&A��k����ȓ(� rs���`��Csf˄|,�P�ȓ&�^ɢ�Ń�~�& �m��%Z��O�!G�$�/t[�;W"пR���
�~�!򄋅a;�p�F6a�
ز"#��D��M�&�5�?7=�Iiq��k@�
*	ZU�7F+>����D��RJˮ�h�`�F]�O:$h��b���y��I'f��p�o]�V�0	�Ӈ��y�ME�V���f\�N�^�I(�HO��$��H��j4%� ��-�ӃV�`�}�������6I󁋅��Nd�`�*|O�7m:}�f�8J�F�Pg-��4a��½�y�<U| �`����|=��K�0�yB�ЍZ4r����v���Q�D�%�y⋚�A���I��@�r� ���@�ў"~Γ_~ ,qc�K�i��Qu㎤XHxq�ȓI~�l�b`K"|>"�!'� y'�M��I�<9��U�tⲍ�!Y�>�(T�Q`�j8�$�rQܑrC�+3#�Aj��CE�5|O�b�H��cџI����@ߤz�j�P��4D��sf�� <�8e���u���Wb`�����8��5k!��1h
�qbƀ7��C�ɲ>Kf� �N���;Ch�9B�	<|����Q�o1�5��D]r4.c��b��'u81���6H�\�{C��=w1��I>Y���m���ɅA9,�˰�X8p��¯G�)vC�ɘ<�J��J�w�L,9�F-B�D#=���T?�8C��'|,RAçv*R�(��0D�Xs#�Q�ca>Y� 5*@AF�0D���qŊ��]�c��$Sh�kEb/D�l�R�QV�����j��y ��+D�|!P�.��a���;�X/(D���NV�QcH�F!X�+1�!�DH0D��pq�W@�n!s+@�&�ȍ�T�9D����iO�i��p���NnN�P*O���Ƽ@�ZՐCn�!Р��"O`��ch�L�.ul�a�A�d"O� I�6�C�4ݫf-�<�p�Y�"O��kv��</e� ѧ�/O�l�r���0����)�^pPvkڨi(����c
` �dOF�t["88'&^�@����\Xysm�`RY�G�wG0Y�ȓqx���A&�<�VPr��=Px�U�ȓ5˱�C�mm�й�d��V�j��6�����iDp�0ebW�Ti��ȓp
�,� ��t%)pF�P/���ȓw��1�`��2qz��Q�G���ȓL�����/( :��d��j	��ȓ�D��f���Q�VD�4��Pb�U�ȓ\f�p�`e��Nt�I��;����%N���	�	����Oĝ
�j��
�1"L-Y�$� +#U=Z��=;�Lԥ�j��a�D^�Xp�,�ȓ�^I�M̷t�2�k��b�Vy�ȓ@����Ք�� ��1̴��5���"�G{�����kń,̰̄�
���Sd	!7, 3����^���3\,щV�J:
�+�L�u �%�ȓE�lz�$F&y��H<�
y�ȓz�m�Q�شq��e�%�Q6���?�nY1Dޥ+�f�%e��Q�,i�ȓ4:���98�X��'��3�
��ȓpZP}�6!'��A�"ި%����c�( I�Ar>����F-b��e��C����Xr�,و��2V.���FP������8�c�k�ԭ�ȓZ��}��L]YO��0�
ǆ8�b	�ȓnUb|ɧ$Q	Zv�Mx���*V��ȓ5���`ņAL�8�mV7`"��ȓR;4�#���]�:�W%C�N��ȓ�|=���Z�w�������*��8�ȓ:@uK�Jw4m@��` ����R\:��.9���J�N[�;.D؆���IZ�S�lqP�!�S�ܹ��,	�}cco�7e�����K,��Ćȓ\Y��{�!�8�� ��¤��e���eH�p���!K��^�=�ȓ�F'E�Lz ��3��?~u�ȓ4����Bϓ�즹I.	1r�
��E�tQ@��,L�`��Ű���ȓV) �;�(J1�ڡ��c�
���`�ⴅXu7�	ǫ�!�V�����{a�+3#XPQQ��<8�X��k���g�x��	�͂u��%�ȓJ]��#H�5'�()B>P�����][gL��^����wē� j���4$���m>0��L�$��W��ȓg���jD�r�S� �1H��ȓ2����ShI�r���:�`ѫt��ȓt�l(XG R�n�X�1���z����ȓ-�;�*O& v�uR��I�0��ȓTg����[�|�4���˴]�\@���"!:�(�8��=#ţ�
[���ȓ$�n���j���hYT'��}��I��Y�����w�^��8S�$��ȓP��"�	�,?�8,�6�� ��S�<��&{�P��#��'}��e\Q�<�Vœ�Y�m� . 	Ux%{0�^F�<هWkj�@����+*�x��C�<Iǌ�����n���&�2d�J�<!Ӊ	PQ<�5�p�S�/H�<� �1I0�QN�J|�S�A�&�YB�"O���Rc�&G�2eʠ
\<A��ٲ"O�
���� �|���(�,��arR"O�лţ�/����a�2f��K�"O�|kV�LAR~�b�T���"�'WR�'���'�"�'^��'�R�'Y a��/�<���X��
����'q"�'AB�'iB�'9��'�b�'<Ѐ'��s�d�� O�8m0a�';��'���'�'�B�'7��',vQY#Lȕ!�M�ϗg5b1at�'�"�'��'`��'���'?��'��H.ľ-�b=Ȓ)ߴ��<4�'���'�2�']��'���'��'��`��)+R{�-b7�l[H�µ�'�b�'���'\"�'mR�'Q��'�h��`�-kd� �-�,v�����'��'���'@��'S��'4b�'���6-�|ȥ��� ������'�b�'Jr�'�R�'zb�'�B�'�x����<!8���[&~
����'�r�'��'�"�'���'b�'ɲ=:�d�9�c�'L��dЊE�'R�'f��'�r�'
��'���'\vS�k�F����t��
��#�'�"�',b�'��'��'��'�b遆A��WFy�hY-wpՒ�'��'�R�'�"�'A��'z�w	4q�0曘�@� �	Y�~��C��'��'���'���'+b"��>Q��'ް��b��<U"٧�ۍ�IB�-�OT"�R�J����$2�d��<��U��P�����;{*~���,*0����M��N�$�|��?	�ѵ7i$jv�¦�VDҥ&D��?ѓ扏b��uJ�l�w^���;a�֌Vźs���z���I
a�|Q3�n47�49ґ��2�n�$h�\3���#J�ve�'���=P�	�je��ȟ$DV�;��L�w�n܁ �OT�b����>>@`�xΛ�w��m0�@�77�Ȱ��%T��rD�'HR�j�����TH~u�˟P�1Roc�! �@��}RƂ�	*�eQf.��t�c�(a��n�O����Quyr2O�(rS��:]`��F�$�.A����Q`�H��_�Ĳ<�I>)�c�;p0l��<a���.������n���(���?A1��b~B �>A���?I���7�B A��*���7D�����W9H�(��a�<!��i�"�$AZ%p*v�)������'�z�����
FJ���`\�T�䭺ӄI�H�
�'t��D�@xn-����'y�	�p,JuI��M�Ԅ��8R��Ƀ�Tup��:?!�i��\��O2��Q�
:��"���
p 䡑#C
�{�(���'	x���!���̾�I��M/m�U��d����Sha��crH�)Y��}:d^�`x��gP���6��?���?Y�'z��u�*R�W�-P�%j��H"&��$ǜJG�+���O��d�O��I�%f�i�O���!ƽ�j1��o�� ��(2�hp}R�'��E�~�K�>�`h�Oo@(r��'�Z�I�+T�D#u
Bӛ6*J(z�󤊘H[�c�'�0���Y�����3�fH��F��z��H8U���(:�� mn渄�	�ZL���@���<Q!�םb��dt�A:]^�q��&b��#�4�?)T��W~���>)��?��V&&�N8� _- 0עK] �T�rCE=i�^� �
��<�ElB,�F�}�4[�K�|R��w��-�@�o=���͸�
���H��HZ��'��'��D�X�F��y�
 �z� �+�`�!A���8Ŧ��8���������f��'D6�'�T1r�'ن\� ��M�p��D�0�$��m��~B@�*�ب���|2'�)�u��\;/�[�|J���yFd�9��N�F�ՉU�y�o� :��?)��v"��?��&�*�& ,&�����I��9���?�(O��c���h�d�O���򟘕I ��L ����]]�a�e�v/�Ɏ��d�O�������W�l��q�O�\�[�iZ�m�e���~%
�cA�ת�.�z�.ٴ"L|(9�������d��d֩��d�#��� D#1"A0�+�������I?v��X��bC����i>��	�̖'p�8��,�I��9+O�7z�A0@eY'1/��I��'�BuӪ�DX&\[�	���D�OL𐡏�|2��F��_������OL��'��H(8ٕ��U��ĵf��^wNb���<A  �$1�i�T���AJt�CnW̟\P�:�H0�����?	��?��'W*؃)��Y�Ǉ�D�Ɛ:�N���A�C�p0*�O
���O����E���OFDmz���`ED&S*�CGCʒȹq5���d��9t�H�Iw�@�JT�?Y�v�����͘C�{���C*��m��z���ʝ'82��ÀB�<��KW����Pß���!�/5~q���6ڙ��胳b׶p:0dE/'~��Iޟ�����H�'*d�pwF�#Y�2�'�Bg�%[�Լ���֬0���0IV4Tv�������d}��'�b I�~�eA-%REc���|N\|a��P�5��H@	K�<�7K�@xƨ�t�ܧ.n��O��9��w��pі�4;�2�j�	U�hS���F�OA����O�Ć�Һ�
��*�	�O��d�O�H���**@�3#J�2\�P@%��O�L\�2!���6�'w�8�O�O;42��E�����B/���0�����N���:PH<��wkq��ju���<�v��@��]>�|�r�a-V����w���C<(5���W ��	��?i��_��8+���?	����*�#G�qӤM@:4�ԩ��JH�Vas(Ov�����"r(���O"��ퟜ-��<!%��G�8kt�3(�ʨ��*#�Iӟ@� ��$��8��4�ʟ�Ih�eW�^@H���(� a"��
�n����=j�/=�����^��-��_����6�F���톨!��$a;�r} �e
��"��?���?�����DL�-��X	0��O��m��p�l*�o�m���A�5Od�lZП�Z��#?��Q���	��D���j��D≠�&.{��|��gV#>��h0u��� M��Zw|�9�fd�M�$+��� ���%
�@�2��#)h�����+�"l(ĉ�O,��O���ƥ}�|����0Z�,�D��@Dʙ�e��1���D�O"�d�iކ���:�����˦��IO9��I�զ ZA �U*v���mw���k��M|?����C,!�i>�3��غ��M��yBJپ)��8�T�@�{�|���hO�Z����L�<�!MC
��D���L3�д=��h��ɟ��I���9
����4$R�eS>T����	���'��s)�q�r�'���O�,pCdJ�.q~=��=Π��4ĭ��$IR}2�'��]s?i�	T�m���	
��}Ap% m��]#!�!B���n�.[~�ц��=;Ql��\���'���"��<���4 ��a"���(�>	KĀ).�r�
�N�)J3�'#�O���'���gFҟL�&uba���\k5p6J��!C�I��<)��i��إ��$PC}�'9��ˠ��b���"�ɏS�����'�<q�/\�8�tE�ヘ��y2L�g���;]ۨ���i�H���]9~��P`�
}ڼ5pŊ�O$����UE4���ӟ�������p�O�D���d�'2�ԑ�QD�!�4Ԑ���3l0H@���'Gr�'����>��d�'Hv6=�L�GΖ�e�$��e�Թ"GR�h���O��DC�M�ė#:r�P�Ο�Y[�w�)��3�i{䃎�g>����� 1�x�0O��
l���y�Q��剏�?����FXp$Q�z_�X���)��$�6k]�U:t�	��?1��?�-O�b��hr����O��	6uGm@b�ӣ�P�j����$HW�I���$�O��I/�~�gQ���m�%���^6е���O��)��kR�<��[�&�a���-RT܁�OR
����q�%�!�ǃpR�@� D�o�h$2�苺\D
�D�O����fb��{�m.�I�O��$�O��� �6�z��a���0\�����ORA�2lʕy|\˓+̛&�'�T���O���)��H>D.P���lP��c���Հ���Fy\��1�}�a�S`��<q�[�$e���)�(��W#ӗ�E��
kB�RD+��V (�+OR�	���P�GN��X��ٟ����Xb�qS��UCBɎ�#аq��Tyb�̏C*`ͣ��'V��'���N��I�o~���r�^9u�� � ��D��OJ��O�e@R�O<�4eO����T�u�PУjؿ����a��:��p��qӸ�Rf�l��K�%ȓ��,G!��_NR��9'��ѱ�(2:�� `X�T_�(��#Y�ivB�'��''U� iw�ҟiD��I h��g$ܭ�Fe�0�٧	? �I��M�����D�'��듭?�����7�R>��0hԑ�L!�PcϻG�xH��O�t&������'�v��C%
B�������ʌ8<�m��언�0��%ί?� �����?��?���(Kv��L~�;��y��V3xXT�ѬV7U"� �)Ox���8<N�E� �?��ڴ�?�B���<�V,O�$��PH�B��;�:���b̄i�T�����K�L����ӗZjt�;&�|%��'�d4��J��,a�T!L�?�<l��GI�Hu����4x��8,O���	'�U�%�V����Iԟ�2��03�p1�q���Z�8y)3��Ꟍ��wy�`I$p��Ic�'���']��!ߦd����#�Šm=&�߱���c���$�L}��'��E��~҉F@� �̧7l� �
""���9�F�Ry2�rc��~����4F:p�����n��<�d�'���&���Be??��HC,��'[*��S.4��럈�i>	�	����'�0��iɶ>S򩛴h\�at<�j�N^Et$Z�'���g����C�:�������O�Z㣍"1�v@a�EA�y&$h�)�O�(� P /B$�a3�U�"�󄌨zhDyZ�M÷'޺�y�S�����{�ɕ�E��?ɲ�'��"�T���'���O:jL!�^>��c��N�r� �A�8,�%�B�P<&��Ͱ�'͟���П��S�'W����4�����V���tT
Ď0j[����?	��D���Bt�[sN,Z�(6�ug�J!+>.��q��� ��M�2} �P�`7Oj}
�/L"�y�dJ�-���?�Dd�<)f�d��%�H��T��<s0�E������?���?�+O�m�Ǖ/�F��O*�$GDC�x�a](�\p:T�NKp��Y�"�	�����O���'
���M� s��O�~ � �wnP���\`�d�y" �}Kt��@H�+�^�H,�
l���'�\;v�C֐M�E
¶Z��ň�-��z6���̟h�	�(���"�R�˟���ڟ�A ��in�`.�����jV	Kٟ��+H:�|�	ퟴKٴ�?Y��NA~�wQ���Gr�jA����pވ�Ņ�L�b�#�'�z0"wd�a���:ẅ�<"��ipc��H�t���Cw!�W(�iӷk�5�#^�\��V��db ���?	��?��!L���(@����
P��ଌ�����=�:� �%�O����O��)Ӝ6�5#��{�*�	}nhСZ���r'P�h�I۟�xwm��i1�[������i 0g� �-�D�f��䀐! y�E�7�e�8����/N2��*�ʓY���K�rܠr�? �1�Eł3JZx�KäF(]���'r�'"[��QZ�?��,��I�}	@��/vu ����Nv0�	4�M���j�z��'Tꓪ?��'��Mcc
7V3NU��؍Q~4����	�1zɇ��
��d3���5�f���iV��i��� "��]�O�~E��6�J�o���5&�������$���qV'?睬SuF��r�A�B��!��'4�������8��%'��s�&r>��I �M3��c��(͓7�e�I�@�4 �	S@�l�~R�{�8y��uC�����#w��<;N,�%'�-��.�
1s�h�U��T�i��s��!A���&������'~�'�,@��\ ���E �Z���'�R�$���P*�R��Iɟ@���?Q�sd��x;�b�C'����V�u�"�:��IџP���C���=$�T��7�Ĥ�Q��:,�/�Xp$B�I%&�CHA�
7B�'���Bܲ��?��`��O��"�HyRA��;���
�G�mTJ`�sÞ[��$�`�D�i$�'�h��f� �I����� '&���*K�� �6\��B�4�?��AS~�"�>��v��u�2��7 ��O��k��i��*c���!��r���<�b)��=֝�"2�(d8O� T����|�:dJ  j�1�A�'����W%H���K���O��$�O���L>; r˧%�(q�!ܴP�>��V�\r4-���{,"���?y�����
[���LŦ��<�Zt��-(l�*6��	7���Iן��R᩟�ǪM��'T5�;4�Xs�'�K�B�/e���ȳϟ�G2e̓J:���5�o�0��IEly��O��2Uo�|����>��AE	�K������m��$�O���ɶD���A]Fi��������?�#(�Qp�)e��6�p`#���?����<���9���П���#��>?�Z�b-nxHU-s:����)�d	�'����!��9�04�c��<yZwna ���f���}RF�{��W�OϲшS�Zx�D�O>�Dx%p�3�%�i�O0��O(������Z�Rd�⣎�7&2����a`��,��ٕ'6��O��������"�x� ���>��$(s��BR,Jg�B1?���I�2{�B7�Fܺ�q��1�y �`
}�;㈕�*кV����$@� E6J�9�Obpʓ
����1-e<�RC�'���'O��Gҗ[(L���!�5Q:��iG��!C)n�X�P��iGŊ�)�
��	ß\�	�?j�.�5k��=��F�3y�$rrb�mQ�	՟���*��,7	�pqʟd()��;{!��B&R�e`���� Q���w� �D&�dPM'X� �{����&Q�`{�)�����'��n��X	�R��F*;H����?!���?������ڈ)�P�����O�l2`�Q0X~��aeݬ4pq(Q?O�oZ͟��S�>?1\������ٴeȖA/|��!K;,���[�H�i����t���4Jt��v�A,�i����X>E��;X+,�W�ցEϖX�2YRE� �$O�zA$A��?9���%o̥���c�*6�H]�!_�GL��'��1�?���?�&Ǝ4Cp�b,Od�l��츂i�@��b�,{t1O$�4k$̓$[r�I�c/���P��O�I�7Vb��z����I#�̐�kN�IS�����6A��l����^�}tl�'����r��M�ā�O��O� y����� �4�Ix�0�[���O4���<Y�,��g#�����?)���
2�ֱ}�x)���)t��q(϶Y��'l^ꓹ?��'����SDIH�1�I �CN�j�J�"w��`�hHrM�1y9�IQ�k��p��AS�7O�dl��?!ɔ95{�I�x�����Xx�<��� y�p�:�.R	2Gk�?���|���?!/OD���y�릌V�6qF͒�L����h��Oj�D��e�	��L�W��	ܟ��w#����0�I�'d�& O�ҟ���N�Ne.� Em%�牼-K�T Ĺ�����yM�*2��H�\+#�r��E���?�d�'~Z�r_m���I�0�I�?-rQNUQ��
Q�PY���O �(�d�æ���J"Ȧd���'�R�O��*�^������k�b>4�N�!��	?�b�Qf�ƀ�?A�rp��<7~�DD?J%�]��uWT*6�ٔnP�.'�Eyā�?t�x���?O�����y��Ǐv��ɉ�?i��	I�e��j1p���
4V���1�!���?Y���?a(O��k B�,�<���O��D��HUPAwI�9e蚑�Y"��dĳ_�	��d�O������DD&J�;�@��>���`�ǽZ����"�P�y2i�f{ܤsǵi����Y>�H�}�`��O�7
�.� � �-1j���E��x֭���?���j��eb
0�䧝?��Ӽ3��̌Wa0�OT 
�R��m�$�?��Ę�N�(O�hm����a�0?�;L^�K�K�3EN�)W������CR�#H�Y:��pu��� )Β�u7D��d�Ea`��Zw^�� �n� �<t�ŝg3`�x$�H�b.�'����V
��]S!�OR���OL����H�*)@��6�ع�&�WRL��d�<��S�v��(��?Y�����i����[�R��:F+��O�Ԅ� �D��i�O��D�OXd`��O�4`� A���	��6��b��| l���/Y�P��&�)�r��<O�I2�f9�?�W>^�ɤ�?y�@�'ֹ�p��;$D|9r��n��1����?����?I���?1)O�#�"�V������=�(����;z�&
�Dߖ*�������5���f/�����ߟ���3)ڦi�!VK�X�K��:r̜���U�&�����<;�z�)f�Z9��6�	N9哔�K�K�w�H�@�^w��E�W��)q�j�s�l��?a���?Y�'S�SL~�;fj\jg)	�\!��[�nJ8gv�8{)Oj�D�0KpȔ�!0�����������$�I4&�L%����7`f,�U-���dc�弟L��L�
 ��4���B-n�A��I�<�榙�R��@A�O�A�,q���S��ar���O��Ժ����haR�Р!r� �������+���w#�~���"���؉����h�'{:Q��">���'p��O���-
3J�fXy�*S�)
5h����S}2�'��kF<�~��D ך�'���r�F�����N�0���y��, �P��iS�(9g9O�t�@ �y����K?�	�28ِ�k��ԔQ���e���-��D �ҥ�?��|���?I/O���;W:�i
�!Ŭ4�4=(��]��B$Βgy�h�8�_� �	����O��8��2�\��7h�4\����+��Lʆ��M6��"���y��H�l��᯻z��Ap���MރNͦ��%Ɍ�z'Ev��O(�	�{@�������h�	ҟ�S�|�rїO1F� ���qh��G\����'��(? Db��'��'8�4A�����'i�7=�����C?He�5i��Ն7�6����O���]+����!)�ϟ��5Iuݡ��%PK��)��5�5���G0���ϓsm��h1.�Oj���G�~yb��Oz��G��q�n���L�Fi�`�E�0�h�C���#��D�O>���Orʓh�����e]$�?����?�%�G�I����@���`pP8%���?I�'Ko~Bb�>I���?I��m?�`�ϗApVd�U샸wy!�l��P��q.r��Մ�9&��/?��X�VZ>�Q�C�O2��R*Kt�萌Y.^�>�i!��^��$���?��W��͉�MS��'�?����?Q��j$���ߦ�6�Qr�۝�?ɒ��-k���)O\!oZןp���*?ͻ��A�6L8=1��D�r��y��4B���'Y��ϕ�u��ɒmw��Inb��Z�M	� X�C/%X��ԫ,RT��׬�剐�?�$eV���B��?Q���*@�P�ZL(��N�Ӧ���ȍ*] ��/O��;�d�f̬��O���X�9���<�v�������C�,��-�t�\,,���ן��	��D���R�J�jG�?	� *���\�i7�	�����Q� ���`���Xd扊7�t��'�P���<i��'���Ӆ)F�iB�q�s�S�[�:Ez �ʇ#�����'���'���'S�	�YX� 6�X�4��UǒEJ�d�� ��4��� Rܴ�?��(\y~B`�>����?�1 �I��hH ]�������Ʀ�J���-��i�a,� �D
�T�M�]�M��a�7������e��݀&���`L� )�2藚>$dhሇߟ8�I�T�Ӑu�4�%?� �*�sԆS�91�R�d�a���������?bJp�Z�'�@y�Bj����[�f���;B�w� aS��K�$2�^�S�O�0�����"�O_,����`mu�����B+���b��T�<�SȀ"]��P��?Of�P��<y$�'�^�K�"�<>�r�'%rn����`���3��[DO�2��'���)v.p �	���T��ܟ��S<iC��:��	K��h���+��Ifh,?I�T���Iş������p��ܦ=~�I[�"��dzVǡ=�P����"��]��K��n��K�	���OC�����=/���Oxy�%kC�Ngj��d��)r�N⟤�2ǅ:H����I���Ο��	Iy���[��4f�pY�������L��d�ɻ;g�	!�Mc��$i���' ^��?� �N���!;D	�����~b�1m��������h�2�p��r��*�`TŜ��y"l̫&1PXS�����.Ыg��?�U�'l���	�mb��'&B�O����S>!b!� {��Ee��5�A���6��a�S����	�� �S!` �SߟP����3w$ҶQvCJ�AZ���$[(�?������)+"X0$?f��9�uw���\���#���:Qk8lY3fWI`�)t2OPGi���y�+_;r����?����|8 ��m���J�.X�~����|4�����?���?�.O���'C����O,��$���豂W�h��(Sv
�j@��Q��	�����O���2��O�k�H�y��	�%��K�K�c���bS�U6�y"���tz��4�i��P�Q>Y���p��T�"V�0��V��EB�8� �+�Ƥ����?��=����ƴ�䧕?��Ӽ3��	:�6A3��юL�x ۃ	��?q���zX�,OD�m�ɟ<;�9?�;`pd�갍���&C@�C���f��"j^���'V<H��h�޺q��y�@���;87���w�3H| ���	�s�JuâΚ)U�D�Yq�E�p����y�O��M+�C� p2}�Gb$>��,���N%C�:fH�<������D{��jI1�|�㆚�mh���\� )���?i�^�R��^0� �2	%
�)��1Ze���a��M��W�Cw��c�eМj�ϓ��T'�O}�Ysy�c�O<}!��H d,~����t|��E�
�(N�ۤ�'m<�r�@ز@"V�tCf ;P������5�4�y�Lb�H�dϜ5������d�O��,_R���M*p�0��}�`�ѐ�����:�-�7W��D z#Yw���a'�k�dn�������k_�U����̨����P�ԃ��O����O8��87����NU�P]���)g��l��hB�7���$�OH��C�Լ !�?�8�4�?�m��<Yf��j�t�k0$؜ZV�����æec�'ld���+�~Zw[��v���Q�3,z�(
�F�>��UbEP�|EP�b�Ř�
�4p��'�*�s�<)��'(�\�bK*���'	�#I������ų~��D��(B�'g�I3y��p���������\�S;��13p,P�y�G��%;h=J��&?	�R�<�	ӟ4�AF��;�L��d��I��^zҖ�#
2MH���+$8����\"=�l�cS+SJ��<�S!u7��d»w=j��'zГ�nD�n-���@�Kk�,�1"�O"\��A;�����O�	�O���<����%<�^��P Pz�z ��m&�m���$�?�������'�����O6a�'�«ԥN����M�x��	 c���ϋO\����"l���K�'����M׺o�,P`d��-1Ł�Z�8M����8W�	��?Q�kK�}�Ƚ����?��Җ�H.���:-����߅i&2ӯ��;�� j��M4���O����9��<	���y�MG)^�8P�oƧ['ֹ��ݱbZ��Oz����ⰊP�5jC�Х�u7d�"�|�K�m0)�l����R�8G8�r�>O��#���?�ï�;Di�	5�?��T+*Π�q�+���(�d\K���OŷQ������?a���?�-OL�QW'�$�n���O���}̍A��,>�Ib�͝.���dD�a�����d�O0�I2�~��҉j�,9RE��7$Z����#�&�xhh���<I2�|�< ���8�i���	�5.S�Q��݉���m��d{ ֶtQ̘����ɟ�I�؉!k��L�%?���ɟ��I�?�FЂT�[)d�l��gF��w�R4��:_��0�ש�XyR�k���䆾6��iޝ�7�Ҕ@�Ĭ+b�Q7���A��)mM~y�E.��4q����<�;	|�b�'O���'����h_j�m0&��6j"1q��S(]d��<q��'z�)R�T:?��'k�O!�yg)O�4��@� ��i�A�O�H��ɤ)W����j�͟�	���?f� �����7C�"-�.���X�*��CQ���$�O�������)0�y0ȟ �@�ò�
�/ܖ0��]�Gō���7mY�dX�;'�V�9'3O����<��'�n�pa�ԄX*2��N h��J�W(j����'g�'�r�'���瘹L�ğܡ�WV(��G2{~�I�ݟ�[ٴ�?y�n]G~�F�>y��~R�O�z�@ w枖^\p�ڱ'�5�q��E�[ Fu)c�i�8�IС{��V�g��Q�-�� ���/����-M�x��@  ���1S��s)�y�	��(�	�?u@6�Z�s�!��#��9�`��6MK<X r���'���Iퟬ�Tj�#@��������4�?ŦI�<ac�-_��	��q|m�"\7�z=��W��xk5�����3k��;� �8�'nഡ� ���ê�&8��݀A�È5����+�*�?�s�	V����?��eʓG�e{��?����Bd�QO����A
'H҂$pr���?�(O4x��H̳>�V���O����6�Jp�لq8zA*fd������j�	b7�ɝ��d�O����!D��A;7ѾC�O��IhG�i�V�#�n�>F����ǝ4a�҇g�=.��\��������ԉׅ��$��[�E�c�*-�ؐid��;P��I�l������Cğ �i>�	�ؔ'�2u��I(��;P���T�aЪ�#ȥ1�X�XY�4�?BZ~"M�>��k�(��#&k�4 $�
&c5���j<քhRi�1�4�4C[�<�F�K�!j��݆;�t�)�3O��/*E�#�V��PP���?!��' ,!*1jD�"�"�'�O��PɀY>�3�m����h�ۧ*9Pc�EN(T)��*dMϟh�������4���@i����D��WE4�ɒ�[)*\�śǐ �?q�'� �	��Y`0�?��N��#�HM�V�&��Ŋ-�Z\3��#<첛' �t U�����$����d���z��Ob��I=_+��0�G.c.�4���x�k����I�0��Fy���_�֭���'��'jVYҶܸi� @�B�A�đ��'-$��OX�'m��'�(�B�'ǆ�����e�c�M 5,٨10��6xR�ϓ&,XP�IK�M�����iŧHY�K�B�;w��(�P��ܟ!�<�1�k����ğ��f�_���&?���؟��ɟ1�2��Wh��k�H�іN#>�����h�DLBs��ߟ4��>�M���i:�E�y7kD�W(�eˣ���`0&�2��+ �|YR�ܽ
�c�i��TY���RT��g���ea�7��inM#6f�?DI�UBB&W ,���*\��ɦ�?ye��[4&p���?i���*4m�pg��.Yf����L��z��@-O>
⪚�EK
�$�O�����bi���<��D�9\�p�O [��:���/��	����ɰ7"��	�s�6�"��?���k�7t��H�� �7��(p��M�2��L@	�n��	�I �#3�'��e�3��<y��'��ek�YS�du��Ǵ���,�@�W����?����?!��?�,O �G�ݿBʜ��E�Om�U`�mÿ8>p�����&\^�$ͦ}�I�o��n�I�0��J��
�&�>a�%X2�ٍm��<��GUm��G��-��̂`L�"]wA�Ց��o�4+��u�AKއw;�a���03Rv[BI�~�q��i�OP���O����4"�ؓ��n�O�⽸�B�LJv�÷�8f^���O:���6E���<���Dɦ��ɯMb�	�>��{�cHA�h�3�mEHF6m`?�-��E��Ӻˁ����u'ˍ�s��z��6*5�z��b�!��?�?�R*�=]�	��?1t���$ H��?��2�xd@���S��P�a��\����?�-O"�:�  9�ʓ�?1�'	�d��C�T"?���cU�Q�d�f,�`�@A~���>���~"���ҁeW�7��ԗ�`�⣧�{�R�@P�O(g�H�y*U�/T�Q�g�Ouq��O_@]���{h|"�Z���'�j[l}�$hR�(����?	qED>bf����?�'�?����sZ&Ȉr�]`Ɋ��vȖ]�aE��Z[��Lm���'�.d��O80�'$�'4eM8��8����x����"��ܩ�+9X��}�pΉ�<!r��9��}���A��g�h	AL�aܤ�� #�$�8�[F��O�����e��]rk� ��ԟ���c�(��O�Z�C'�E�fwQ#Q�H:+e�=�am��'=P��'�'���'���a�1w�I��M�;f��r>�6�Z�&A!�
h`��?�@�N?q�c[;
	v�'��И\w�`�f�2^��0�wi��.�s�䅣%��Di5�)r�d��0��nyr��O|-S���A���I�وG�̷,�\*d���]���OV���Ofʓ}�i�b���?����?I��RBU���)QF|0�1��?!o�W~K�>!��~�㡟�y�ϋ�Iq�蓡*�6����޶c��r�6O���ț�O%Dlfi�� ��ӜjX4���U����W�I\l��I�Y��j#,���?���?��(�)��K~���?��C�I�ԇ�UNT���;~(e���fS�T�ǫ����ئ=�	�	���Ӽ��J�4�4� �D��\�ұ �Ӆ8F�A
Î8�?�U��8��U]w��I�c=O`�ʀn �u�
N�6����I(8�L8����*f�a��^\y��OP�qg�͟A�����Oj�$��H��!`ۊL7*K���-,f�{b��Oʖ˓o�^��#��?y��?!��e�v��'�?q��I-��i 䋓$��0���/��I۟��	�|���� �4+��?9�a�w�!�f��M�*��5�����nZ)�3�z��@`�̫ႎky� �O�<dCV�,���"��;$���ҵ�ʄ'�:���O��d�O&�D�O��D���y��R4�?A�B��'� %��@�<]_� l�&�?&�ir�(����d}r�'��D͕8ö}ٱ!�zaV���!�9<���KQw��ͳ@'P�<��L�=���]�|��dPWQ>	���aa�1���=]"���1O�8�	9vt�����?A����������##	V�8���b�KJ�B���MR����O�U
"�� ��:�M��+�T͓���OK�d�3�#P��KÅl����{�d`e�^?�;C�<dy\wV��:O��8�e��D7�����I�1�^3��a��om���\�$	� s�T94�ǵ�?��?���8m��r��ҧJn
!f��
���O2˓KVRqf��?���?a��fQ� J��M�(ā�eAQ_}�̀���M~��>����?���]?1#���N֬�S*F�,�5d��Sn����K <f��ϒ��d8!\7�6�����'bPZ���<��� �`���>GEz����׫Y�Ş�[m���`�'h�Ox��'剄H�̹ڧ-�"\�eK��( �[�IV' �hM�	�����4�?��l�]~ã>��HH�!P��N���TO�nq����A����ڧ#���q!̚�<TƖ<ɍ�;ml�6b�#��5L�2�2�#-PD@s��O�]�ɚ!�H� ��������������O���0���-�$�8v�@�" �AoݟG�"��@�'V"�'���`�)���SȦ�%I�P��+�$�b��7	8O�X���hb����Pw�OE��$b�
�;c���� z����"9�$ESdꚶN�"ˑ2Oh��2g��y��%
Y�	��?G��H\dHc��4#�x���ل)��5⡉��&��c���?����?i+O�;)���#��'h�'�(T{�D�#��[�E8q����'ZJ��O�E�'�"�'�\XJ�'i�⎢!����ϙp�(YA�T29Z���a7O���u!�� G�$�CN��:���\���D�% ��KtiM$`f�0�#��>IdF��ƅ�?���?��
W#�L~��?ͻAw�qz4�(j4V(z�A
�ȭx�l���S�(�?q��V���'"��O�Ԍ?@Vy�P܈v@�<���S"Z@Q�u"M?+@��ʃ��Bh�3��<�b�D�`�}�,��w�'RL�5y���G,�x	��ּK�ʓ���"���b��'`��'s�4��&4d:��B��6\��53q
՝tL�
�T�P3F@=z'B��Iҟ��	�?1��]y�g���e󡇘�� �(���t��?��@q,�Y�"ѩ��6J�G������M%�L�␂B�u��ݱ��>ي	ϓw@�O���3F�[y҃�O �Ɂ�9!������d��h�2݉W����BM�O��D�O����Of˓<���8cEJ�?1��_�ɐ���	0�����?��i�b'����D�G}b�'�R�Y#eӸ�� $�W�؀[�A�	�P�3@��,#�����.�y���,Ǽ��;s::Ÿ��|��wb̢�а7��A����M��Q�
�vP��E�'=��'C�d�Ԝa���yg�.a��U�@<E�=c��XgUR�'~�$�#3*r�J`U��+�4�?ɵ���<����6	��2�.��rBr8���n:%��0j@�$���ta�;(�Ʃ��'���&�`�*p�d�RYl6h��.��Ol`=ϓ~���/O����!G@dX"�@ҟ���ҟ�A�����.�3����)��uA��H͟���my��� ��0�'���'[��^-I���C�'Z�z����^�YM�2�O�p�'���O����w� ٥l>�z��^��򐊕M��4�JtEY�yL��	t�ǞX�PjV�e��	��~ς X�Ҫ]�-�gB׷@6E3�J��;���eʑ.m�b����H;}��)R�ZF�D�r֭�� s��sH���t���Ϛ4Y���8`Ã.V�$1s��	����H�!�+"������#�=�>�3������@c�J��84�B��0D
�6B�.� �{ �7�F��'�w\\�����y�	������дG�8$��X:�&�--��ak�ͷ���cd�'�dY�-96֨���[")j~��A˔0/����#�(M`����#'���2��� �|���i+"L8�*�:*�HZU*X5v���9�O�-��:O���H7���O�R�'���1�-J:[������}~:�*��Y(��'N"�'��\���r�L���Ǉ#�`��ǈ*?n�\���7�M{p,��<Y�zd8��?e��ʟ�1��>a�@%4��!(J!%���yw�m}�'O��'��	6g�`�2��:��@�z�����fe�s�g� �֤)t�i|R���~���?���=h
�b�{ҁ��5�쌀��
9j��5���M���?I)O� 'BZ���'zB�O���9�IL*r�H��h�+�"�s6���~r�
'�?���)�5Ex�|�Y��	|�.ujd��}(�q{e�v�Vʓ
��9���?y���?1�'��D�N���Za/B#������ {ǐ��6��O ��N v����4�dX���Od�e� �1j�!��I]	[�4%y��A�i@��'���O`��LMX]�4ɠ�
�0*y�=��!C�&���z��i| '���>�1���d)]~X��Lȉ%�4]�D,� g2 nZ����Hh��V���dH( F�d�O��!��i͚A�E5ɊAa��T\���}�c��_��'`��'�"� 9ض�ʙ����U<*�D7��O�
D��<���:�?���v���?��3]
"��acV
��Y5���oP�L�U����D�O�d�Ox˓G�����,Xp?�U����w"�!�J��~!6N�Or���>���O���'I6���G��8TT+e珯;�ҥ�WĘ�/}�'���'O�W���6�Q����`��0�e���cc���U���ҟh��7L۔�韒�d�O
4�vJ����O�g�q�!f̒u�P�u,�>!���?����$&'0��'�?᧡���	��g�z��D��t����'�Dؚ�'9�LA���?y�N��'��H#i�'d���X���hH;�4�?A����$-��%>����?ט	��t�:)�fR"_� )�Y��'F��"�[���[w"����9O�n�6fx�����-�$����˛�\�4	A��M��\?����?q*O(���ω�&�4�P��؃%È�	�S�P������Iݟ��<��MC�BłcϜ�k�.[� �l\��D�ߦ��#;�M����?����"0^���9�V,@%��q���!��r�kăJĦ���G�ڟ���A�)��?���7q;���4n����m��yX�V�'���'>�-�a�<���s>��	�E��6Mǉ|�)!&�[�J���FY�&�'#�'
��g~�_>7-��'KbY�Ƭל+��t�'�H�Il���'z���cU�$��{>��I �韜,1B(S+zs�e�")W��B��Y≷q�P��?����?�.O��c+]�?����!D1YI@E� ��]h�'�����? �|��<��`�q0�K��b�l#4,KP��l��$����~y��'�E��ԟ�u�f�ͨFJ��c3�Iip$;a�i�p$j��'-�\(�~�'�?a)���Y!�i�X��7��$VRy	�GB�)��ExK<������OP�`�|Z�p����fJV^���9$��70z�IP��i���@��~����?�,����xBˀ�%������-g�~]���MC���?�-O��R�՟d�s��Kq�݀j\~���g"4��ʐ�~"B�2��dF˺[���?��yZw��l+�Bu�|��W��+ ��yq�4��A��lZ����O���@yb�ȹZ�R-���Ġb��P���5�u����?9V���?	��|�/O���� �E��n�3n�Q�C�@��L�ǽiD�����'K��'�"�O��	 Q���,t.t��e�tT��⨐�VS�X#�'�*���!�Ş�?��V�.m�����0yX*|3#���n���'��'�@9�q��<)%gf>��I��uh�� ��X�k�T����]��M���?+O����d�O��d	��{�'D6B�̭��B�� �lZ���+���dY���'�P8uQ>�'oH!x��M"⧀G������&�M;,O���!���O��<Q�_>~�*)xTf�H�f�AҀ�$o�6Р`_��ÂM�O<��-p��RyZw9v�ʅW:�F�]�n�N8�۴�?�)O ���O��d�<y�H�	S|�)O�(4��K#%6���5���~�bo
$�?��X-H��S�V>E��]�yF꘻;Q�Tp�M�7X�j�x�O��$�O$���<�⌖�~�Om�eI�)��w�D���#-���qӾ�$]./r� �(A�i>Y�I��'4���R� ��k~�<+�`� Y�]n�H�IUy"��!7j�����k̊0Tre�!� �Km��RFD�!g�`��vH�X�'-ם�l�)�Ӻ[� !u\�s�b,�M�.�z}��'< <Ps�'%R�'��O���/9_�3��8M��M���¼����6�V���ϓ"��0��e'�S�S���g�WLD� _�d1�7�(U�~�lZҟd�	̟��ӑ��D0R��Q�K�(�B��Ƥ=�Z�A_�RL�0lZl������ �1���D� |o�Se���NfT)��إ.Œ�o��4��̟P떈M����X����OD���i�.���^<zڼ���W�V�ܴ��jx!�S�d�'!��'k��Sw!K$VͮPP&���3rڑ���m�,�d�(Z	���'�
�ۜ'�����yB��5ց��|&��3l�1�Lc��Đ�M���.�"�̓�?	��?����?�.O(�b,�?���I
�C�vD�"��$)���'�ʔ���?Q����<��'�?��Ut�JE 	'�B,���q�⩁��-}��'���'��T��!m��$��5>�<���N�xC%,���M��@H�<A��k����Z���?9F��<��8'\=�g�C�,^������`a�'WB�'�[��I�E���)�O^=Ra퀧sزı஄�]A"��cHɦ������	$@���ٟ�sjw�L�O��+&��{�� ��bU�sn�2f�i���'v剡t9H�������O>����yDmp�mȀq٘�%��cZjK3O������O����@(�(��F��ci˶C��tX�M:M%���r,��i�'�P	���;v�'R2�'4�F�>�҉ՖM�<�S�lHs��
`Y7������?q���<aK>)��}�S
Bh�ve�)EC��h`�N)OU�7�D<#�!n�x�	՟l�����B9^��Dn}}���� Vz1��F�F�N(oZ�=!��I�ؔ'�^�I����'�^�@��N�q�^@1��[b��;��w����O���ƲB+@��'�*0H�'T2���M�uʑ�m���3CeM�/,�LuA��5��Py�ȗ��yʟ����O��䑎!:����ĀL��;��Q�xnǟ@T"�*��Ĉ0	e�$�Op���4O����.\�$�tM�<H���^����Y�(i�g'�����	��'N8 
���bÁ�� ph�q�φ���y�$���?��(R�<����?9�h��4����]{8E"3��990��i̓�?Y��?�-O\�Ɗ�|bC�1Vyz@�A��,/e�]�A/�æٻ�e�t�I������?��	ן�7�>�aX�D�թ�A�(uҼ�j�jO��	�I��Iӟ�'���#�!�~���{Q��$.�"�9�MA�FU��HbH�ŦU���#B�扵M�z�	埤*z�@�i>7�<�\��@��
����h�X���''BQ�HD�����O��d����rJڽN9��	F �NJ&m��)F��]S� �D�O�`C��H�'2��w�ѳ���p�)�L��F�7��O��\,o�dmZ��x��ޟ��S�?A�ɺW���z���hm�@c�,���q7-o�(�IJ����'��	�\���Ӻ�jܺS�L��d� )7�`iA��ߦ����M;��?���2�W��b�n�l[W̊>l� �(\���!1M�0�M��@T�<�/Of�$�$�1����$
�2���$A<��š��zļ�oퟜ��ǟ\I������;;���Oj�Á�i��qpui�)O��I�7�պN9.��޴���O�m�3=O����l����tp�MJ�2�� s�)�ljt|��G��M��D��]�� Mb���ɫX���	�?��+)TY�bD�z�|��$e�(���,�r�����O��$�O����h�&)�ڽC!�_(M@t�k��Tb�	��\�	�삳�q�����4��-�X���`{� ��`7�j\���?Q���?I�����ۻf4�8�'F�<��t��u�湲wJ�xlZ�lZ�5<��D�UDg�P���L�����5{L@"�J�t��tJ@ �g��alɟL�Iן���yy"O
��<��?)� /6 �Cn܏�bJc�6-���'b��ѝ'hb ۱�' BK�y��>	7�+^�b�+T��
�@��������˟D�'�&p���5���O����J�V�q����������[6\8e�O,����'��$�y��|��y�1�B9Bφ�B�l�:%
<�bex�@ʓ[̲x�g�iy���?I���I�X��8m�2<�mQc/N?\x�dc���O��$����)�D�(c��O�4qB"Z�A�*d�D�8m��L ޴I���i��'��OO�T 0H�I'Y�T�B�+|$��y�KT�6�޴&��y����*bDy�|
��2b��a��E%qvT��瘣|C
�Q�i���'�"���#���4�*U����b��t�܋�.ڪ9|����n�s2���i̞�O����O��F{�? �X�Ǎ	�5�eB�m�0�Ǹi�BN�2C��ʓ����I�T*!�2��%��	wM�"{�hp!�	�k:���'���V�';���	���'���ƃ�z�@��E!�������R�f��˓r���IʟPÕ�-Z��?y�h��{��Y׬�A(Q�$�����ϓ����O����O�˓|k��F8�ƐQ�K�(��o� ��D�'�z]���?y��q?����T�I5.+���+]-�\�ǧ��!w��I�#	��èO���Or�D�<q��
)UA�O�]x��Vp!@�B#�Ǝ����+vӺ��~S�� \���'R��R�'��rL�!���ې�������n��T�IryB��N��^���l�)��� �]�f����`�qRF� ��D<��'@PI��'��'�>�]�J�tq�̓�t��\�3���UH�6-�<�%�ٶg�&G�~����FV���3B�6�F��Ff�#6�����OZ�	�<Or�Oj�(@��T���	�!җG�	���׷�M{� �6X���'���'��$�<�C����A�VK���EKç=�F1�e-U��M�F����?�L>i��ȩ�?���*�0;Fo�Fjbӛ��'���'�<�(��<Q&�k���ɿF�7�9�d!c���b��[���#�ObzW�(�d�O���O�H&�4l�����_)8n��Yw�U¦��I�gR0-O�Y��'�r�T�����"�3�k�[���@I��!1���C^����n^ǟ�'A"�'%BT��r��	������wu�  "��l8��(O�q��'B��"��)�O����W��2'b��nt\��Gk�</�l��fd�O���?i���?�/O������|�
H,w�*�k̌/{:;�\���wD�O��*A��O�b�'*�1�f�'Ab%�4�ߠY�]��M�ň��@J�>���?�����:N �%>I����d��"���=3'Ԅ�riD�M˜'�(�_u�	f��'v��*}#��	�/V�mA�I��^-�n�⟔�I��I�5�]��ӟ ����S�o�H��"Ɲf;�ׇ0Y�v� 4������O���꺓���s��u'��
-"Bƾz2u�`'u�ʓ&��!��i]R�'�?Q�'��ɍW3���S��	}"�{P�HH��i����1c��HZvC!�fglQ��lQ)oɸi�&�#��$Ȗ!�"�'�2�'���]��[��y>1:C B�JU�e" I�k�xu���?�Q+��}o�#<�|b��3B��4#��i��E��#�0բ��i�B�'�gL��c����Iǟp)qe}�
��kK>>���X!�I �xm�Ď�;�1O����OP��ڮ�V��GlC2sT}�$-ݪU�nʟDj�&���Κn*�'B��x͟k��kw�-Ô��	��� �S���Ajc�|��ӟ �Iǟ���-m6�iҳ#�qYj��F(B%Hg��by�
�C�B�'�&4������y���UZA�%��@���Re�d��&O������O��$�Ob˓���9���'��2"�d��g*d��);5�i�腊Q�'}�ܕ�������@�	><�5�j��v�ٛ�GM&s����?q���?���?�fo�<�?���?���wp6)q��`�f�/�Z���i�����~R�'�?y��ґg�P��Z
�Y�A(G�.��`���ˑo���A&�[��h���͛"����Є��HY�,��3"�!�D}�*���öy��z�C��b���L�,$.\�qGX/;�x���q��b c�>
[�%R��ǅ	�2A�&@(�h9�Y1�V����O,{�ɪ�%��M�hu� �:E"�b�曫t@
�xDT��� �D&S�i�F��07�R̉�#V�xZ1�5H�G^��8�C�bJ��S��a����A�����Ob���O���q���\@E�թ��s8�w�ZT����<j����'HC=�Ƣ��~G�g�I\l�r�A�E�Ĝ:���F�������g���b��4�$/9�3�d%��˃�\)�z�e O���O��3��a�i>�G{��ٻ_޼{�a�ct������y���� _<��懗j�.�K�kH��M�=O$����Iiy"+�"= �pu$��)����10�v��+��W��'���'q�4�a�֘A=b:��A�A��=Q�`bm�1��$  �܂��`4&� �!Q0�"<OFܳ7̛ *h�����&Kь@�bB�	�b��s`@&{����+$<Ol�CWeS�5v�`rO�qQ`$���ur�'�ў�?�Ǯ*l��a�6���X�Em9��=ѱ�$ɱ!�2�Ӈ
ؕ4e����2K1Oz�*�3O�ʓh�����<��'������A��/S�Y������?���I83������)�p�: Ap)W0c�2ak�i���c�=% 4XE
Y����	Ǔ}0y3f�2W�����M��M�cQ�s�I�ՆV�
 tآ�j�8��yW��ON�Ĵ<�v�C�;�jqP��<��.�|���=��.R�BΡ#:X�C]�nz���n��y����o����d�BlVm���<9.O:3Q/ .c�
���O��'^FI��`M�'�S	n�H7�ǻr�ɪ���?q�e���C��<� E��O}����g�(�O{��q��ŢT�@0;Q���R_2�J���ed�>c�r�H`�� `	���)�*� �s�n\9a@�Ʀ��Z�s���I��M���?9O~2���T�(6�ࠡ�ћ+,~�����?	��?q
�C�|��
�8Kz@)�E�h�Ez�q� �"/1�S�? BP����r˰,h�!��ha@���'M]�D9�O��y��",}i��ٰgY=�"Ox���%Q'?\�1R`K�NV�C"O�fƄ�?�R!�O��iK�0af"O&*�7U��� mS�K�Tx��"O}�7�4n	�Pk�
6�,�"Ox��N]:e(�(��Y+iZɐ�"Ot!���C��}�k��+�̥�"O�h1��s{���E$!r���"O��"j�gȔ%8�Lĭ���v"O^����8+�`Y�K���E;"Or��n�B����Պ��-aP�(�"O�D8��*'v4���jӻL`h�r�"Ol1��eּkfJ|�JX�	Tl�B"OZZ��+_����Þ�E�t�5"O��A�"O�O]N�(WM�*$*P� "O^�85*OJL:A��

�,�G"O�e�D'?o�=:�
�]�d�90"O��b����^ PÉ�x���@�"OF�2�k�0\���Q2{ؔ%:�"ObՒ���'��=�1��-��5 "Oȝ�a)�]�R����"1"�ʆ"O���HƚWw���a��A4����"O�a�F�b֥x�\�$@|�3�"O\�86��/��lq�
�n#�A�"O�!01o��"f�H�u	"O��@�"O=Δ�ԧ��qy�ը�"O���4Gdi8tf�$WQ�=��"O&(���=H*<�e��=;4���T"OL ��%�������L�><��"O.i��H��lp�w$�12��q"Oإ;a�]P�@��%C�,�@��"O� �3m�,���.���S�(D�D�V��
m�B`�پw����)D�cr� �_UN�HUa�w�1rK"D��ȑk�<X��`���ɫ?�d���>D���6h��Rn4���N,Z:h����=D�ܠ6��C�V0�@b� ��<D���Sށ����� rI8�@?D��qtFI�0����fiO�gE)�v�0D�LBp�W��e�0��95���IE�;D�tI�,������G�!���yuD>D����+ЋLCF�)���W1m���=D��k����x����`.4�&�;D����DԞ�<}I'Ɲtȝ�/D��`�폜F�|�u�-�T�x'F.D��YsJ %O��� �"Z2�,D�s�f
�]�c+�D~�1@'D���C@Z#�����(�p5b?D��+'^M|���!s{��#?D���%Q��d�Pg��a�$ �d!<D���B� ����&�na��I�%D�<�QoR(i���.2���j$D��:�%8-t�,sJS��M��b#D�4��
 ,'�iBi[�ol�y�@c3D�h���"3�m�P��'%5�1q�0D��x"�܃k޼P�tBXNq��`l.D���2)7i�N�%�{6��`��-D��(�*[$}�,�!�!�Ccd�B�h-D��`�N� Hi$�jCn�ALVV8r!�d[�-tD`e��F40$d\?[!򄂧jC���&�o�~a�e��!�D��I��*E�����E�!�4>���a�GW�`��!5�k#>C�)� �����42P��o�t�1[@"O�<k*X�!��8s��ˎj�)c%"O�{fiY��l##�
!L�I�"O� 1���=��s#]<S46�0"O� �EWQ,�ӡ؜?2��3�"OѲ���ZP����AF_��I�c"OX ��Ñ�7O�`R3@۸4�ք �"O�Hh���s�&���b1�"O�5�@V�z�����N�1"�@x"�|bN��Oq��+�lF\�r��S��	r�5�"Oz`���/5&�)�-N�xW�h�`�xҊZ�������9�3?	F�X�z;QQ%i�a��T����u�����+ 5��>�@ݍO�%��b��2��rR�q������牋-�0t�'���I�L����'�`�AaZfhiF�G�$�"i��n
Hmگ|ɶD�	�w`D8�(W�E���ci���| �L��'
r�' v��@��
��� E8#�,�9�hF���i
�V�4S� ž*.�\�ƃ�q�ɼ.&�\���\9��Yd-^1�B��
:?�o�5%*q�c$�b�
D�c�G V��]�U���?)��P�|�l% g�U2��#�	�mzN�F-�_A�9�%+\A�Qۢ�đ+TB��L�:��SК��lZ�|J�O�u�� ��@eD=v��T8dNL�L�p@��T�$�a�EE�+���$C*���JO L�MB�̀y~b�'�����>�D�(��S�K��p�3��'�܄�6ִ?qj�?��/^-��d��p�BD�3O](3�Ê}���`��8?6�(�&
�}��4*���|��3x�6�*�.�=q��c�>0��#b2�
QҦaڬ$��K�H}҈�4	Sf$�-#ĉ�G����h�'�,d(�/�H���/�W<Xq@T�|�'�5�XpBP�R�B�X�Ն�̸'Ӣ=�7�H�=g|,rR��G���2%���;�k��B  t�wy���%?�x������F�3kD*?�V\��ǈ	_��H�dT(q3�O�iTJyb��=K� ��J�3�� 	%D�A^.�/O��dN�Qwڜ��kW�N;͒�G�#_b�����طD��I�]fȖ'#�cA�0q0R}zT㑽48|t��V[x�|xP끝t�|u��F;f���"@6/⨩�	�4Z}�e�ec/Oh�j��vy�*��
��<����1���Y�%]9`j�Tq4�XT�I ��Us0�H4H8́��]�%��➈�s��6�Ţ�JXn�ra��(��!����	ӓ|Y��-G$D!�ɸ��r�Z��ď��iYrE@�������0��$ҫ*�jtxZP�B��p���O*�ِʏ=P�����[힕C�1�I�'eйj_������-��dS
mdx�0	 �i>����ϡ�$iϓ)�>����߁^s$h�N�7ORx!K%�#chA03�O,Q�*]J'�����81D$�(O�8p5�$�'= ��1%�zL�7��ƭ�M>�3�6PƬ����hnQ���D�f�<:�#]�Y@R�XS��Rd�3<O�+��5`|"T���=�LQ2#[�.]�/R�| �,ҏ�O	MS6;��dhD��  ��=n�>{]T$př|�'$�ų��w��uY ުkU���dŪu
��h�&��Tx����"!p�I�<�H(f�	����RAd-cţ^]x������d,a��N=Qt���/T�YC�K1�؉!>�\���zB��1l��T3���+�Uy��I:u��#7�PH �UT�.$� �E0.�U�Z2Ӛ���0�I�&�Ms���&*	������OW ��hOQ>U@���Kh1�UΞ%O�.h�&�C%^��c���e�X�P�T>]��E��K�nÔ|��,��KE6�5J`�J�I��4Hh�j�S�4M�b���K�yKf+F��i�1Of)B��-)��#��J8����\�dΓh��3������PaX�$�򙋲�
O���iG/pF��4�X2y�iD�z]�Abj�_�^��wȒ)X�F��ӭa&����=�IW�'�`�D�̉�:X��GH��X��'�ȝ�%�'�zu�� ��pa��O��h�=I�5%N��*b�8hj�����DGA��ڲI.D˓.�L@�ʍ/L�i�7�ɩL<H����1+������&?3�P�`o�x�r�w&��p-Y�A
N�ѳ�`��dJMW�d��Tz8����I��
��Ӥ�!cu$�1�4�I=M�x-c!.J�gjI)dB^�>�ԓ���p�S/J.ɨ��4J�*8#
e�<��z5`Q�V'Y�7�n4Y��(C p�K>Y���,K�?]3�w�&Au�L�E��!D�K��'vƅ'e����p��}?@�xbgL�uZfX���-����h�����1V�����U�d�� 1¬PJa|ҧ�uv�;�8��pb_	.0�P;���L�d(��_��#�P�"j�(+˔�%����p�[a�;F��#����w @��S�? � �b%�:Np`m��EaR"O�M���&kbX�[�'u���"O�ՠ����~���@ϣ)x^Ix�"O<!��c	��x ӌ��{a���S"O` DNНb��гī�%SIr��"O�4ZU�->��[eϩ-&v��"O��u�@�Mn�����+�Lu"O��7��	SҀ�A hF �@0"OL`(��@�p�@̢�F��}+g�?D����$�/N�ȑ���2Vp+�,#D�D��Ƀq��]��b;ؤ��r<D���W�q_HYC&�"صBf%D����& 5����媇�.d���8D��pģP�x�Lq
�����Dd�c�;D�\#�S@1� ��F%�Lp���$D��A `V!@�𻁀J�2���$"D��	Bf��a"���H>D��="�G:D���ԟ+Jι*Ee�,u�Ӥ=�O��	�CM�r��a!e�޹e; �҂G��l2�SD�ҽ�yR)~�v8W
<d���@�V��(Opu��)z�f,x���T�ibi�`ଂ�k��DFPL�ȓ0�0���/�|=:@�҅h��q
3
B�%! �B��a���O��Bb�ӏP��Ah�=J��`s"O�mSj	%�\��rܝ|QF]8T�O(�d*T�g����
��Hhh�`��b��Q⅔Y�48���	-�`I0B�	����g�Nj�x9�̀ �$9
�'��)8��δ
��Y�0C�&3N1�	�'T����"8���B\�	�'P��i�F	�*�E!�V"�)�	�'�\`���P6(� $��+�|$3
�'���'ᒐfY&谇h�2|b��'L�h��h*<%���]�!3�'�Lx�IRb1�x��
G�i"��	�'�,�ddďr��`��܌{�\�	�'�L���Y�mdn�	u�z6)
	�'�8�ZW*�'|�j�NϙG�d�y�'W��J��vE����?x���'�m����9J�<�jB
�yB�Y9l�Z��8l�X�p��&�yBj�� �̵Ѱ�30�� ����y�Ě�Jp��ΌY��=�����yr���3�|��#o�TV����nV��y��V�e���:S#HJ؆U�2J���PyA,�$��-���YQ�<q�ġ����������L�<�6�Ba�A
�M�D�B�ᣧMF�<� kD:ꈔ��
h@:�ɕ��h�<�6�,�����ɑ�6�%�2Fh�<q��֡8��y��X��>�hÄSy�<�$�տ�^�R�h#����s�<a��=M=���B/ �4���1���p�<)Q�bx����8��4�эx�<Y6�S)8��)kVB_�#��]�
^[�<!��B�n=
9�a��<:�e���l�<���ĖwȈr���4��`�i�g�<�3G��Z��tz�G̲SDx�'�@g�<�d�ժ_w�:�$ɘ5W���ǌN�<i�D��{ri���Zj�n�gJ�<1⥓�%��}�MR;�Er��OB�<���� �wΙo���R��U�<Q&@�/F�B��ֈ�7X�l��e�F�<� ́�$X��BU
Ԯ/�(ӄV}�<��f��t��uCO(� cfQ�<a�R0 �f $�;���Mx�<� Z)���I��i�Ҩ�j���"O�$d߇X~x���@��v����"O�ehbY�.��H���0=��쳠"O��h�'�z�梌=*��X�a"O�h"*ܞ�Peb�B�?}|Y�c"OT�V�H>b0`�h��k`6�# "O��L�X��栔22E~�Z�"O�p��,�/l��*�,0u"O`c/F$L��"	���k�"O�xȇ�%M���B�#i� �B�"O�0��7�D�`J K�!��"O�tp'��<�X\���-�� "O��:��U�Pcu�2��J�l�x"O� `�h�*cݒI	4�^O�"iA�"O�Ҁ�+4��
�͛o�ja��"O䕩�jˠ[����@M�����E"O�Y��.�H��qP��#kp�p�"O��;SF�#�|C��˚?�"OX�9�D̟2~�iZ0J&]ײ��"O�=	�G�Y:�EI"k��bZ�Q"OtX�C;\v�I���OΉ33"OZ�zw��g��!��4��$�"Of��f��L�I��֣8���"O��z� 
P��_9D.ށС"Oy�'"D:5��s#(�,<�I�"OB�jd�����	�8.�q"O��b`+��W����S���bM��"OHɢ�C+<��+���"Қ��!"O��h_�QF����H�ܺ��%"O��)s ̕K��p�!&�����Q�"O��"�B:A5��k'�ϟ<���q"O�4Z���^�&)�c��2�@��"Ofѣ����6��t;�a3l*	��"O�c��ϭ~R�$ѓ�R#=��T �"O��!�$Q:yJ4z)�#@�Z�:v"O�����0	I�GCE_���e"O�`���Mخ�Bw�!b�Z �"Ovpҵ@]�`���ˁ�S0ۊ�qG"O�= ��5�8yJ�Kf��i��"O0�sR�
 �f�Xj6Dy���t"O�h��	G�I�8��(�Xp�8[�"O��1��gW�^���p�"O,�c7�6g&:w H�^����g"O53� ��\�*��F�v{~쪆"O�P6�Y� Ѓ��&Ml��E"O���n���4��\g~���%"O������s��+W�X��0H�%�y�.��N�m��~��ز ��yL�
h\���J��X�)�n���y��V��tp���(U@��w��1�y��CVH$�b�ƼvX�)���yr��/B�,�zE� �|�&�֕�y�ɋ�[����V0z!��2cB��y�n��|��؟t�b����	�y"�L�y� !c��\q���;C��=�y�f�J�Z�m˫[�"-�r�@��y2��
90j��E�NА���y�AUpY$��b:@�f���K�y� 2���f��aJ �y��A�e]�Y�hW;bXD��QKҠ�y�G˴�c*�S2z�҇N��yBc p`j�R��®O�A�-^�yr�ǣ)F6� 4�M�Cg����.�0�y�@U#}�����A==�,[r���y
� z��`R62�ʌ�6D��wA���"O�i� �S	"X��-ɶՔ�Ѱ"O��R ]m#�)���S�4��y+�"O�8�"-��8 �,�{4�8��"O�	I0�	e���#�؁W�$��"O�y��"�^�x͈�O�+��!"On}�7ܼ���r���+k���P"OL��4,��K*���N�	��M;p"O4E�`���&(B��29H�4��.?D�x��KD	L�|�d�&y�����7D�,���"����悖bK���&�:D�ܳ�o�TJB�r��N�Vڬȴ�.D��&#X0)�|+�+�BFv*��-D�Ƞ�	:�^9��
�@��D8D�P�+�
��ȓ6��P\]���)D�HS�H,3f�j��ĵ']���V=D�4��iӳ0���k�%D�q,��I��>D���+�_`A�
���j%�)!D�����.�`8��H;v�j@���4D��S����b�R�RF.t�7D� +�G5rz���L�O�^]ɑ@6D��R��~�0�x�lh�I{�!3D���R#��E�8t23�ܥG�Z@p�1D��H���rz�	�MY�w� @1�L1D��#Pm��_h���X�k���):D��AP�R�n��$�.#:��@�8D���V\D7��C��'X,��2/!D����� �6,B�JѫvO6���� D��І���7��p3���@����� D������Bh�aT�	;LP	��*D���v�\?��ʍn��s�K�B�I*ܬ$��]�Co�`��l����B�I�x����WC�:~<"�ȍ'��B䉪88Vd�S�B!2�
	 H���pB䉞A��	Ӗ�Ƴ���af�
B�,f��Zeo����e�C�!���^��+럷5��aP唒z�!�	�\|��5a\��b��1�Q6H�!�D�/�*H��&�Е���+�!�G9>05;`&�%�"\��e��y�!�$�r&B<�6c �NXP�ˈw�!�D�8>����\�jo`�)5$	*tJ!��D�����h�)�̾7B!�dH3#� �R��7�@���Dݥg+!�d��GM����~��pB޾2�!��Q�q���[f�0��K&!�$?M���j��zDp��R�_X!�䘕C1J0Y��9yҜ�k )�l�!�Ĝ�]�:H�#�"q�k�-޳s
!�dP?S�E�W&�-'> 0�LK�r)!�� vt�A��<=�����/�!��0T.ДX`(��e&8���o�>�!��Dv
���O&�XM��-͉uy!�V3t�ZY@v�ׇZ��-{OQ1s!��:C5�:$@Ԟs�y����'n�!�Dx�f\Ad�)��An��q��I}��H�����1B<�BR�[8g���2�"OX��a�Os�X!AnւZIr"O^I�%��2%����l�P
���A"O� ��蒬a/��0��6@�IQ"O l�Q�S�v�!��*S37ےP"�"O��9��+����z��(�"O��{��"��ɡ�B߂�<�c�"O����N�"&�'Ø�4�0�R"O� R!6���<�~H�ퟤm֠�w"Of�q,�РX���j/�D��9O��=E����0x�h�"LW �a1"W��yb`+[��L"s�KP�萮�.�y]�j��4�h�G>p��0�/�y"���P��Vș�	a���u���yK�v��5X��Y����e'=�y�'�>r@�Ұ���O�,a���
�'��[�D 4�j���D��� 
�'�daP`��A6�e:,�<�:	�'m���b�Km�DI�*;Y\đ[�'
�K3�ٱ4��(���XGFD{ۓ��'��
S��OlXU��"
*i�;
�'	���S�/l:`�� ��
CB��	�'��Q d ����B���-�8:�'�����*"jp%hgDِr�� P�'��}zգ  �P��lD�����'�t�st�kB b�n�Bx-A�'v`y�fS;9�e/�iR��
�'+^l�WKXkʍs���<'�t:
�'���9��'0�T"S)�t�08��'�pT��K�<��dh2��	�.���'����!@���-����	�'���jV"� ^�L�3��t9�'����II�.��9eGP�'m��'�.����I���hQ�̀6�LXJ�'�ļ�� e���"b��9xM<�9�'�ha{!��^�:5�� 7~kX���'�B��&Gć ��#�i��A�"�!�'Y$��At���(ױ,3�w�<)f��<y�+&�=%BB���N	v�<r3��T�2�� ̪2��W�<a�.ДВE���Tņ)2* V�<9c�ِO�t���������&��|�<�&@S	���(&�Z�S�X��`{�<I�ҏ<t�+�l��X���7�s�<A�G�]��(q6)��޼���q�<9�� w��dk��i�˗��g�<@iS��6���D�m�B0���c�<�&�N����i�Ւ���G&�Y�<a��L7��b떏B QX��{�<9�-ʏdް����CƜ��#J{�<����%i���Q'G��]��w�<�ҢG!�\�t"z �@k�m_v�<A�!���$c�D�x�P4��q�<�Ri����{0,Z�Y1,1+$@�j�<��m��+X��0� �3J��� b�i�<ـ����jЦ�-��d�
�~�<�č*"�p�� ��D�⑳r��`�<9�H�R�H� ʁt�0k�ev�<�a�N�&�{�fԻm��k�/W�<)��ƽ3N�aE6��:7�Q�<��̋w�&P[qmƲe�)ҕ��t�<�㤕�C��Ƞ�҆l�J "r�[q�<!� $,��APe�� �.$�+	W�<����~	�D2���9 Z�X���[�<�d����zDj�,n^񺗯9P_!�	 /nt�BĒ�H�@�!�mA�]!�D��@�����3����%@M!��B�����j� �r$��DH!�Dػ@�V��dm��2d��xD�\ ?!��X�����1��p�ݩ'��$�!�$V���X�J^�~�N�V�~p!�2^��e���um�5��[�!�� h}���X1@��@��FM�)����"O֠�q�#yU�I�G�(N���"O���G�]y@2�I �(M2"O qj�D'�\h0"gЋ �.��`"O4�#�m(<(�����T�Ju"O��&M@>m�ix��Z&S���r�"O���$�U�37Z��p�ls��[�"O�P"�G "������K�tБ"O��Ab�o#�L���ɰ1��xa"O�I�ㆧKh(�6� $6Q�"O^!�B ��uT��i�L 
i��s"Ot9��������,a	Ơ�""Oj�3%�}O4�SK��΂�"Oh�;a ۴3+�T�#J��S�`��"O��Z���Nh:�	D�D�H2"O1�3��+Iz0A��
������"O��[Ǭe�e�f��:]��т"OV0:��+j�����?cl<p�"O�������Bն]��啾}e�-q&"O���d@G��D�'��s'�Qx2"O,m�"�Ȝ���娋(Pv:��"O���E�%ب�VjXI��̓�"ODbq�U�X�� +gh[zJ�d""O���C�^*&y8�t-�*J�T��"O��8��X��(���S=�(j�"O��;�B�?-��*��.$��:E"O�����@:�xv�OotJ,	�"O�W��c�#T�I8c��d0�"O�]�T#W7-�ڈ�JD����"O���$f���J(cr�2
���"O�	�%X�^l6]�0��^@Ct"O��Qꑖm����4(e9%"O>YQD�S	���W�.�`��""O�Ѥ�E�JF���ɡ�v���"O��x`��>EJ�����Q��Yz�"O<�Z��3A� �+�%��+��aq�"O�)P��$b�eց̋�@-�f"Or�I�k���A� D�|��c�"O�M��������m��c>�S&"O�P��J��{6lLuN���"Ob]��&GR]�P[��43��d"OJݙ��Y3
1J�k�Ν}/艁�"ODU3�-�I+:,���ÒVx��"Ob�ʲA�r?P4��E�	c��i�"OJ��D�M�BhH�В�Φ�8T"Op�g���!c�<Y���SR"OxɶLK;3�Fug�׮��Ep`"O
0a�'�3A�lQ�%Vu^̠"O�dC󂘵4�j�a��#e�*�+F"O���� [�r�lHK�Ń�c��y"Ojlr��Ѕ� ����6L�F��"O��2��9[ 
x�g	:p�n��"O<,�Ѡ��4�-V�D&lS,�C�*O����Q�"�<�xT [�&	ބ;
�'Ŵ-K���n���.��"X��z�'�,����P_�J&`ɼ1r���'�X�HiƁ���+a���"����'�1C� V�	��,�q�")����'2����Aq�S�BJ�@e�	�'F~�갪��S)��cWI�;�n���'�v𹐯5��6�hX4�#"O p��C��209�Z�x��B"O����IN�t�M���j��T #"O�X�FJE	jd|Q�5�K+=@�"O� H0yw��W섹�fT�6z;�"Oz��(6�RA�׏��V��{4"OH$I�ަV���Κ+�` ;�"OjX ��V�{��8qW.�Gx�) "O8��T!\�L	+�͘�zLa$"O��c�u���� �ؑ�u"O���k���RC.��6	���C"O�y30`��H�Ơ����?7ڌ��"O�К�����xUf�)��	 "Ob@�ge�=��j���"Z�:�"O���a�,h�x�Ze��n�֭�d"OF�B���)	��dc@�$�yd"O�i1"яR�P����,z`!�"O�Z0�׷nM"hK#�#`����"O�qĬ��W=�u�$� YȤi�"OlD�d-Mr(�SR�q�(���"O��[@k��O^1R�� �I��@2"O��E�3JOzQ���Z�"�3"Oz!a�'�3;8�ye��y���s@"O,�K��J�X~H�U`E�_�*D��"O��!ߛ!T`���� �l���"O�p&(C����m���"Ol��`C_�	��p_)|V�s�G�<��N�?ŶXҗ�^�f�h�dE�C�<��	ֱ��㥤��Y��t d�C�<)V�9:����BP�jM���Y�<���\�{�Z��.ژ:Ͱ���JU�<A�˔�!ˆ�����Bt!�P�Q�<	�M�UF��M�<K��X
0*!��)�u��J��&0�=ab��v!�$'�$�D%V�}z�mG�9�!�YVZ���וpn�K��)�!��J�#�4�� ��CX������A�!�$���X���g�wT@y�ʌ�X!��Z	C��8$#Ϝ'KT	���M�u�!��"���)C4=���@��b3!�DXpH�``�Q�G(:�+s��-3!�DYW���i�u:3��2;/!�R
b����Ł(�X���+!���.G�>!r�G��4�x��07!�Ĕjd"�7�L)j�T�r�E���!�D۱b܀��6d��A�V9գ_�F�!�d��I�#L��bn�+p���I�!򄊫���E���ȒPl�!��[5R(�,K�fZ�g:��3�iF6}!�$ܝi ����T)t����]�!�Dˊj���5o߶ `�5�!��vΨ�QF��)�Бâ�q�!�ؔ�Ey��ȑ/������2v!�d�YZ%b�Ö�
�S$ᙘ6!�$�6m"Db�CO�X~�H�q���/�!򄛞xLHȐmYha	G�H$u�!򄑆rc��*��N�I����ޘq�!��&+�j�`�K;,z�`��@U�!�D��Ni6mS���.h,�����8j!�$��R>��ZsK��p"�Y�3- I�!��:a/�	�������K�X!�?������(A/Ne��Js!�7��Z5C )6�t�`스>�!��	~�`3g�҆%�D�
E��2'!�č1V������q��-Y /\"!�d���V��W'@�F�Rp���Y�$!��GIpD�4���2��t G#F�!�
�
].���jT>H�N\K��ïw!�� �8��0Y��j�=,dH��"O�[vh<P��Q����NjE�d!�S�	y\�[���W���Q��"!򤋲A��5���.�X����'�a|��R�v�=.&2٫ABK3/�h���'5��0!�ΨK5��Y[
. �4�'	P��'�ٜ2��nF=t"��`�'�j���S�:��Q�J�m���'�@��gYM��1��	w�P���$'�Lࠅ䎃W\`MPD�R�p��ȓ|����e|�z�k��;�(�%����u>�|�d�f�,e��@~��B�I)�T8������'��wD�B�Iy�v�P��=n��-*�AޢLjhB��-ڲ(±A��0���y�nB䉪"�΅�u!W G�^U��dA7J &�=Y�N�Mh��21p\ ��Aϳ#�v,�ȓD��U�3��76�b��5:*lՇȓm��պ҃�fʜUyhM[H�?a��0|BK���/�ȫ�aK����ȓ8Pq�*~9RD��4i�l��O�&aI��@�P�ܱ�L�?m}��ȓ�J�e��[G�h"A2<�ȓB&昣�@��a��Qw-���Щ��0ȺA
Ð>\�pc�
�.;C�E��e�0" )S��}I5��g�P��G;6yM�j �qp���P���1
䨥̞YF�-�G鐍VK⥅ȓa g���Oc�T�B�[�C��<��z�ͱ1�L/<Xԡ&\;,�h%��D{���Xi��ͱO�'3���aς#ў�E{4O,|��瞞\*�2��M,E�rE���D:���D������T=w(D�M��iIў(��I�ц�@�#p*��(o��rT"O���_�1��� l��0px�:�"OX���aG�K�*}ˁɌ>S=\���"O�88W'�#k�	��(@�dɤ���"OBQ�!y�
�#mK>&��Q"O�i��@C9�&�C2E��Y�āx3"O0��������@'��u���"O�A� 쌊<%�f+o���1�"O�|`+\�"��P
�;fP��c�"O�BvL�77�`�0�53&8�"OXP+�!@�G�٩ŪN)}%2-2�"O6h����e��iyujX>��"O6����N5� �����fR|�X�"On�DC2�`[��D�>� b$"O���$���.��DG\� 2��S"O��{R����"�F�6���B�"O���Q�Q�,�8򔨉�?�����"OqC�k�."���qB77���"O����]�N�����W
}<IK�"OL|b��BxB1�T��u�6�*�"Ot0cЄP���SF.�82�0�	�"OT`9B�
�M�8�I�۬F�bU��"O� 5��\	��mQD��x��"O4�"�#j�h  ΢�>J�"O0���-L����ycA�|��R$"Oxy�G
� x4� ��'9�p�K�"O�=���g�ޭ�C�::l����"O. ���F����b��ne50"Od���"3t�'�$G�*�"O�w��1j�ԉ���� s;&��1"O�pFF_�5�ؕB�o��x�"O� ���uP�i�F
e�@$L��H��"On@��m����VF��.jlu�b"O�uiG��6{/Q���q�8�"O�-!nߕ#gҭ�F$���y�b��A��c1�H �0�䓶z�T5Q-=D��Ӏ'S$?1�&'��rU�/:D�t��$ʋ93�,8���B2���GB7D�p���	�Q�*E�o�*���G4D�lC4�8�jآ�
�2���)0�3D��U�E�^�Y*���:��j�I1D��c��U"l"�ʅ�M:s�����+D�\�ĭJ���'e;1��k7k(D����R����zǐB�Pi��*O62+�<e�i��� 8�l�(�"O~a�3�֮a������{�,�V"O��+�l�%?H��	�Վ_x^2"Oݱ0�0O�:�%F<ng^��S"Oh`�e�WM��kv�e|�)�d"O�4�'B5�!0 �T[pB��"OJ�ϋP�`@��Nة%ex=��"Oҽ+ �}�y���q��0@��'��dA��5J��6IqĀ�3F�#4�!�X�8�ԃh^SL\�@��K�!���e�2%;ï�+?�@2��/nP!�DÚA"�y"��ކ=Š���-2!�d b����BRK�8� s�Ɠf!��= k��`נM�{���RG!�D�9|Ih�(H#���à�� 
�!�DI]�$Y1�	�������no!�*AHMC���G�-В�[!��4��]��#,�V8i"��*Li!�#�Ơ���[�	�<���)�!�A�r E	P��8�jyZ���;r!�d� �rtYg�Qj��pq�ďXV!�d�_9�}���O?%b�|�p�Y�j!��
�M����T(A�&}��kőo���)�'J��|Ж`[0,F��C�%A[N�S�'r�m�uC�N��@{��@�7��H���$/O�8uƟ��x����a
���"O �I$^��M�p#[%\�)b�"O٠��8�T�C5��r��R�"Ov�aC�J�]JHW$��E�+�0�y�GC	����S�p}����(���$�<�ӓTAH��T�����)�b��ȓB[j|[4��g:�(R��D���pyU��Od��~�"rŜ�"�.H���1�:�ybJ����nA���M��D��yR=k.�G���.	s���yb�A�d���b���8��E/�yo8:�(��ѧBxfz������y¯6�j<�!�ޙlH����y��4
h�k�"�f	Ra�2o��hO��)J(��K#�[ )��(AĊ���џ�F����%ξ����
����#�cי�yBG�731��OL!#�Pb� J%�y� ;_r�bfD�	�B8�`ܫ�䓿hOq��5��
�G����q�Ҝz�<��5"O| *�&J$iխ�[��B�"O��k���=�As���@���8h��{B�dZR��l݃	Y��)2�H�9�џ�D��W2
ȆP �,*E&H�Ǖ�y�Z�|].�"j�(���#��!�yJ�N: ��#�=���.%�yϊl��܈�-� {2͈�?���v�? .e�GH�	�� JI�DQ"O���ƽ	p���F&�dnAS��	m�O���rV�Ͽ|�冀�%ƕ��'���jP�����!M�N���'	���@G �L�����y6�R
�'��'I�&��t�!��ѹ	�'a�k&�Q�RP �1#���#�QU�<����/fH˦��q.�*#M�G�<����n:����(�i��I��L��?�Óm�5�D���H�Jv�?S��(�ȓFz��ɰ��--8$�qp��!V��ȓ�D\Yw�
3��u����Q� Ї������������@ٽ�z��O<i�.�9
l
�q� ;�4$
0"O��y�cȠg�D�"  ��в "O��│Z9X�H��sN	�:�)UW��'��D��'*Д�\:��a�� �ɒ��hO?]�� \5.��I	�@5H��i���DC�<ip��c��}A���9�,UX��@�<I0K��K�r��D�'�Z]Pzh<��i_���u�N
{@xBK��'jaz�J�b�j%�Um׼"���wh�	�y�C*߬�{�mC��{'��y�й$�*j�c�5�H�(G��(���hOq������I��r�Z�4ޮDx�"O��`�`$���A��7_�\��"OZA4��ݤ�8�f��X企�0"O�i�	K�o�>xqğ:�v�rW�v>��#f�O�z�JFI�� 0T)�@�;D��;V��0F��؇� �E}@M�)�I��|$����~��T�Uލ Q�-�ru��iU��y� ̋76Q3����"�~ 볬���y�O�8�$8G΄�A�P��-Q��y�`
s@�y3#��Hl�xCa��yb-ܴ#TTu�Z�xA�"ۡ]N��ȓ$]l��.F�T�,��	Mpܽ�ȓz�py�2l�u�0�᠂�/�H`���~�A�&W�c�l}	 C�6�<�Gb�2vEq��̖\�HJ$��<��C䉸{+|�����]`j��J<	ΰC�	w��Q" gR��!������=�çt���hwB��&�*$�@d�#� �F{��'H�[�È�y�^A�+�9Ԫ�(�'�����5=������ m��
�'X�9Sԉ�:a7��ELE �c���hO?)jp��+�L�ە���u�:i�Z�<Y7k�����zW(��Z{�azsNW�<Ѵ`�+8��\�4�O#� 4*� Yh�<�Tp�(��AK�r۠xᄍ��'�ax"����@��4<b�i�ƒ�y"	Ѿa�qP�"0�a�U�ȋ�yR���Eu��J6�C-����K��y�gZ�R"���ݮ&��5�D�H3�yR�QQ�|�V�F�t����l@��y�&�B}
=���|Ȩ�a��	��y"�@`��+g)L�n`2L�S#[�yRo�$T�0�GN�w�*�sɜ��y2Ñ�k.^���$O?w��탒�`ɇ�m� �k��x����l@��洅ȓN��#U膂mV����wފA�ȓ=0�(C!Ha�(�q
�&���� �څ�N�Fn���%n�,�ȓRd}@)B+w��)�E
"x%�$D{��O�6�ҁb��L�Z\��b�R��i���� .�"3��9y.��Х G#��=�"O�9�aI�h~4 r-�9uh5x&"O��ѡ��UƶٲS,�;A���Ss"O�b��Q#<���E/��T1A"O$���3�*l����<0�"Oq�S�ٿH�f�9�7��tr��'�ў"~*VH�w��P����@Z�<����y"�y�n�0ī�+t�����y�k��o�D���EP�
Q�aɊ9�yR%�4���{)�sC����ɒ$�y"�P*�`��qY)rf�Y��+	�yroT�:�tU�2m�k�օ��n����?њ'�z�(���7��X�W�F���hO?��a@�s�R	��L�ID����T�<��� �zs]�jA#1�f!��	
\�<�`��2j�̕���˟8`܀��� W�<a�O�!T���ۛ�n���IO�<�'-OG���`��1⌵�s�u�<YE:�T�`�՗:�=���u�<��
�.a�Z����f����g��n��?Ó:^��%j�k�ʽ��J��K�n��V��4	(5��eKA�L����A�>|L>պ��?U�ф�#ݨ]���
^Jܱ�q$@՜���O�p��0��`����ǖtD�4�ȓd�"�o�=l*2!cB�Ka�����j���V� :��,�L�y�ؑ�IA��������,Cʘ��!��o����5D�D� F2�t�H��<v�e�f0D�x�臇q��<�A�O�^#����A:D���b�;|����p�Kn}Ry��m=D��;Q�ß�>���GDM�1�;D�tKea_�k��e�d�^Kʤz7D�4�֠ݡg1^9aa6�t���<��0<�N� 5�x��p	X!�F(�nNj�<qN�
�x���+�.y��|����e�<����
��8f��4�x)��e�<�'�ҁ4l1���GF*�lY���|�<���["��b�?��gds�<!P�Y"j��P�-K���ĈF"�o�<��<QN�m��đ2q6��pjn�<���u8��v�ԤXn� %�C�<�1��%TsG��&j[�	�@�<�fDهu{�i�V���Ye� h���B�I�>�<��8g�,ɢE�)=�C�_���W�I�x��c��� �B�ɴa�`(H��IfA�EG�^M&C�IDG����\����mǫ  VB�ɺL��"@�#�V(Z���:B�I;�z�gD�#�V0C��p�FB�	�5-H F���K�6IuT&B�I$_��p��=o�"�U7mUB�ɉ\v��4nV�y��x�hP�e}�B�	7�,���ߪ<���!�Ϊ+}�B�`�Zi(������oY�2ІC�	�3�$���m
�(�rQZ���x�&B�,g����Ԧ7M8�E��]�.C�	�t� �s�,U
m����,*��B�	�?��9[C@�x�r�bƏڎs�,B�I�	��W�1i6����3F� B�=R�� :V���rjpx�䖵J2DB䉟@D�cs��_������X�k�~B�,[NDbMüjm� 2L�	\6B��7h�p�Tփ-v��#T�Ҭ�RB�)� B�gҏL$�E���I�?{��"OpY+�⎠v���#̖3xȑi "O0\A��T�TjDūF�KV!�"O�9:B��:���fi�t���1"O2QA"j�0\x�d�2t��4�"O �
{��Q��#��%{���t�y�͜C�!�������Z�ybl��I�е[�Ο&B6��0G���y"�@�0��ǥX<?��hj ��yo�l(��/6L�[�HH��y"�~��j樇rh|��Ϝ�y"� �|�dq�	�h����7�y�))+Ƹ�1`D�:���k��y��� ���T(������jþ�y��ˋ^C"AqG �7
[v�f/��y�l	�|��r�X��F105#ȥ�yR�u� ���O֍�d�	У���yr�����w �����@H��y�NN}�L�rb�G�Ro!��y�"[x2�O�����ǌ���y�/�v,�U�1��q2��yB/�	�rE�EJQ�U�.� ����y��r��c0�<2�j�#�=�y��
�*����kP�&l��yB�G�d�8�����2_Qf�:S.ֻ�y��ݴ6X��aJ�D�2I��yb߳W�2a�"��fA���A�Y��y���]R���C�V�]k���0�R��y��UH���w�ަRP�r7F�0�yR/�@�x$[�@-M:�i'�C�y��E�a������=|>��Cf�y�+�2��q�EN�b�<�ߞ�y��6?��1'ǌY`6ݘ7Jֵ�y�a�16; ��)�"J"�c  �	�y�
��7�R%����n��'ꐞ�yB���s��i��Ĉ(;Ђlt/՗�y".E7=(RhP$0xv��#��y�Dү9����ө�&Εc��	�y�F�"�&����R�=6����NV�ybB�&p@'H
�<�<�(A��y2���2�� S$��	E��Y�/�-�y�d߻��(8�,��B%D�3�y�C9�������A�ZE�d4�y2���,�0�$bő>$v-�Ԋ���y+߁q����`+�s��yb
�<job�kPB^�t�8�rg���yr�G�m�Nm�C��Ɖ�e���y�N߃���h���	�x�;�U:�y�/�#��k�ݛo�Ner�e�y�͉�>6��:u�	h <����y�F��M�>Eiu���d�2u��a���y��F�T�0�:��&X)\�Q�=�y�K��[M$aQoěd~��L�&�yҨ�|̾l�L��	���K��O��y��Z�U���ԉVX�2��-�y�i���	�g&��G"IV�B9�yB��[�6��,�!>_B�	�@�#�y2�Գd�ܐ�V`G�:whmV���ybA6S�Jɱ��  ,�sF���y��-Ea�pZF��"V�2<�yrB�?E�pݩ7+��^���&��y�E�,�T���b��\v�e�ǟ�y�ƈhR@���#_E�1%�"�y2��`�H��	nږ ��³�y
� �pd��#q;�t���ѩ:�H["Oј1	Q��x蘥DI�R�D<Ie"O�Y��b >n�x�c��ޱn�E�d"O>T���q�`���m���x�"O�LH��CFd�ac��*{U~�#�"O�d*�D�W�%�B�Ĉt>D��"O�ujp��E�ru��h�G(*�v"OH��o]1���ōѼ�T!:U"O��*Cf�4{lʀa�F��(�4��q"O�� ��C&ir�ԑQ�Q�|}
4C�"OĐ�@,�5T�2����;S}"�7"OT9�g�3~��ukgB۔I�x��"O�i��8k���q"b2L%�"O�ћ���s�(�u���eDPE��"O�:�"E�>���sB��2WC\e2�"Op���0XR�B`��%3h���"O�����ٚgQL`�ю�!j^��"O��8g��%G6��b�͆aAZg"O>�gF
� ����E@�;
l�4ks"OL%Y��΁/�ܫ�/[�g��1�3"O��Bs��F��=��܆I��(K0"O�舓��0��#�+Ɠ,熑A�"O�)��^�UD�АE�G�( u"O4lP`aO�q��Es�M�$H���[�"O��hF�H�<�ra��$R�$�"�"O��2O7Xbd{��L-B���w"O�Ł4/����t�ؔ5���F"O6��F���ulD�1�ёb�� �"O���͍, Pi�ғ)�Hm@�"O�H���&uF �3�ׇ7ú1 �"O�a)V�p\�w��I���b"O�L9�ʋk,�ӀfP4YI�"O�ѣ0��!	P���F	��.DJ6"O�aY����@u�e%_��0��"O�!��ɋ�CL,�4+��x��H��"O<y��&�?���d�T�H���Ґ"O`��A��QrD7�+6����"OJ��eN-@������0|��s�"O�`S�/Y++E�TsP#�N\~���"O*��wEŞU�h
S��bAXP�5"Op�CJț�q1n[#:�y�q"O.<C��?G"�u�h�%�J@�$"Of�Ж��6�Ȁ�b��3]��]cU"O���YY-�H����6�P��A��X�<�� О"�2a!�hH>P�}(�+�j�<aq�W�/�(�PHV��ev�f�<���/�XA	g�?#�-8F"�K���0=�/B��يv�:�59�f�~�<��CB�Y!&`aT�ոk\:�h�[F�<!�a���n�k�
�s}�t��nA�<1t��J���aF\�ba�e�t�<��	��6p4t:�#G>OTdxWh�s�<�ᨇ�w6D����!L��`�g�h�<a�Ƒ��7 �JpYڀ�\�y2i�y�}ӂ}nt���y���6��-a�/m�hta�L��<�S�O�6����[��`[&��7`��R�'W\��"%M�n�0�)�
Q+Wt0Ps�'�V��-���0ԩ�%�1|oPd�
�'R 삵&!)`x�$���i�m��')���,��
F�=룈�V��'�ƅ���6݌��S'���9��'�a�@���;�`6�ݛ�����A��QR���)�����&�y
�  �h�n��.�]Bp�V�E�}�2"O(��Ӂ�(��u2�3U�D8�"O&AX�,�[z,q� ЊO#B(�"O<]ۡ�	�}�5/Шl4�Q3SZ��E{B�&iW���㌍K���"!P��FC�I�!}TɡEAɕ8|��eNY�k,�B�I, �RT1���a��=9�bB�(�.B��Y��)b
˔����-�B�I>���C�6n}�x��&�
B䉬'�-C�2���D^���C�	.`s4@� �O&sRļ�Yb0�c��'�'�az�m��h�\��Djų@Ոt�Q����y�"�37�9�Ó�N�z��!
����4�S�O.����KX�7�\ ��őb����'W0Q��!�1�6�F�4���	�'	ܕH��
^���{��\+�tH+�'�~x�v��!����ҀI�����'������I����26fP��0�T��0�� q��qH&U���"Ob�m�}��"��CE�A"O^P��䑞��)��J޺ 6��y"Or���,I� Yi�À�|HH�R"O~trJ٪1��ܳ��I���8�ę|2�)��c��ͪ(�"
��c/H6X�B�&�^����΁��@�V��,�O�����`��Dkn�2d����L.M�!�~3���eV�6rp�z0�L`m!�D�59����ӊ�\:�
借x�!�L�?+J�c��Q<|R�q��%_,6w!�� ��9�+�M�,j椁��DT	B��)�fx��4Y���8��N>AZ�^,����ƣޠLx3��O�㟬D�7OE
��W.�Z�R�L�?l�i���'}ў"~RX6I���j��M(fP:�"���hO:��$�?OA*+�BԎ]�
�S�!��L7Uk�3B�J2>��t�pNZH6!�d�J�X@���c�h��E�ŉ]*!�D�#jh���V�'��(���.�!�DÉ`�(�*6c�L���B�h8a��y���,y�$���V^h�2W$�#�^�OT�=�}��ř �����l��釭��<)f%ض`^�I;&�6} ��F�e�<)PlG
A���eD��ld�B�UW�<QS G�,((\���/�<���U{�<Q5�U?cXI�u �p�J쳥̔s�<Iq�בm��:�n�#���Dk�s�<���<-+�к�f-�:���HF�<i5A�C���2Ȟ\�Lb.GA�<Qd��H������dN ���|�<��EK�<:	h�EEr�a�aWm�<����.�l���g�8�	���d�C���O��͂��W�e��Bb�	'E8����"����G6$�,�#��N74���"OZC� �&R�Ո�X�4���"O�!ɢ�3�H�)�Ō	rƚ["OR����B~h�q�Ĉ ���v"O$q#��ޫ0�d9Qw-P"V����"O��h�*�,O� wj�/"�by�"O��y�!E��
�)���ww(�{O $��A*yl j�)��`{��ȳ,/D��]����D+k��Iu�O9.!��>�	�AD�fZ8��AR�EY!�D�D]9a���=���aM%�!�d�4~�ޑ3U�R���y��]A�@C�)� $H��M+h"hAbG�П1�v��@"O�-a�&�b(������|{��'���',;TU��)}N���V2t]��?���ɟ�5 �C�i��q��G?I��)�T�������3:��IS����U�	�'V�A��)A�*��ԃ��Z*>�UI�'�R@	d%�jt���w�C.Y�5��'��!��((8<;�I�2~��>�R��(34L)F�^._BR����h~JV  ��P,j�(aY�F���'�ў�O1\�S-B�P�R$+7	�"�\ز�'d�U�TN�Q_��@�EG��xC�'T�	��h�i����΄�z���'��k���.⬓r��,6����'���96#Y"�29I���(�F�#��D�Op�D1§^��I5HF�qlh����W�z����ȓ2W8��O�@öe��Y*L D��N� 8MQ�k�d��E�!���� a>lA$]� ������(0k:D�ȓj�Y��Kʨ��ć�N-���TPL�$�@�*)�4:�-������nǜ3�����m�+3�̈́ȓK{��qF�ݑ(��53r`ѧc��-�ȓ%�pM�!BB(�di"A�ԩA<TA��w]x%��!�? � 5��#��!�v���v���Z�'�9j:0�c��1#�P��$��uyA���HS�8ru�׫Z;X���m�p�*��!<.���V&�5��؄�x�tM�R���5�13Dhޅbm��DLb��U���e���I�$-D��B�L�����50�N��W/D�A6��Z�f\s4"�" ^MC�� D�X�P��&��pA���_��(5�<D��P�͈�D���P$��:1��2�$'D�P�&&ݢ�FӠh�.mH覨$D���AA�0���⧎1C�u�0D�ī�fY+�:uwJ�%Q��y%'0D��{�*T�9*c׊H������"D�,���B�A��H���%�Ԩ�S$"D��I�I
,s���#�7��d{ �:D�Q���MR���	1;f�i�C8D��Ab"��DN r��6\��6D��a%O،6�ތ���I�/~�u*�	)D�8�0�rEi�� 腡aC'D���@�Fa5�� �gwQ���� %D���),�>Ȓw��$IR9˵�-D���S
�d
H�/�%E�A�7D�BP�E�2`�� ⛾k^��jG@#D�X���}�`��g�]⬠"�!D��g�O�/��x*g&�� p9��>D��K�A�F��Zc��==��ڄ�=D�0�FK�v��H���&M)�t{�:D��*��9Z,il -c����#	-D�|���B��{ S�b���q�)D��Ab�:9yL�H�+��X3��&D����JV�4�zq�%ՋUС��($D����d Pbp�1&�62��!z��#D���+��S�d�I�h�?:"1�"D����˞�Q����%Mɚ=> ɒ1$!D��)�H�>]X�ҫwe	{��:D�<��g�@��`E��H��W�5D�8#�דg4���g�ͰWf8�q�5D�(��'�TI��*M��Z��H3D�L˒j���I���]Rı��G,D�� F�[�LY.����4+T�h��i;�"ONEq���"����iM�c��9f"Ob1�Wh�Yk��2�.��a�┩D"Ol�Z�N�
yL�`%�Ѷ�D��"O쌓�
� bH)ՏU��}��"O�51fF�Y������+.e��a"O��8T�W�װ���א)��H	%"O����"��/�N����.)��"O�q�UMw^���U p��j�"O�X
�Cvw��2�/�h 2
�"OH�r!�4�&M�P�Id�dm�@"O�03f�&(��"rA��!*�"O��zR��k����� �0k���aT"Ovݣ��H4[�Jy:u�#T�
#!�	)U:D�b�<x��0xVȉm�!�K&x>��q2��?9�R%jv�J�t�!�D�%�J-%JR
?��(��O.p�!�$��*��b�'rD���.Z�w�!��O'Y����ᖪv\�8��(ղ]!��0v���BȐ�]P�Qe�!���
&a|Y:b�J?,�x�=2/!�d_�/��h[���3�A�w N�v!�ƒC�x-Ä(�5o��a D�ު!�$3��H�6`� 
��!���,���t���M���9�e[�m�!�dȬ+l$$8 EBn�8��U˟�C�!��:}F�%Z�/\�?\F\�6jвF�!�$*UW�"b�ͳ9k�(cF�C	�!���W�I7�(m�P�Y��ߡL�!�9`���u��<��0�q�T�<�!�Y3:v`��@�7C3(�ר�1d���(6$�z�!�,4 �sk�y���=o��U�F�L��b��,�	�y�3X��W��=�B�
'D9�yB��v>���P�.��4�F�C#�yk��YD����"���%�>�y�.��:� �QA�,[zp�J�E��yR��!c?�`a �/T12����yb��{%~��e1MY���'��y�J p^�:Rƀ1z�X)��j��y�ՑC�z-��6?��"�ܧ�y�HXy���@
5�¹"��y"$wIx�IWKF�1aD�B�9�y��g^dh�'.ʆ-��@�
P��y2������Cc_�B���pA��y߳B�e8��ǞGHeR0�y�ԛ]�d	�rO�@�(��Ra�,�y�C�V��8�q�W65l�i��O� �y�-	�'�u�����-�B�����y����6���Ү%0�3A)O��y��Әw��qAB&=)��蹠�F��y�,Y�U (`$�[��(�# -N�y�"�s��=�%�ޥ ɬ���B��$wL����ĥ2�$� ��GXC�	�/=��2��3 �YC �&>�rC�ɋy~ES`'�q2VGS+f�&C�1N!H���m*h0�u��� �HC��j�J0k��C�U�r�B�-��B�ɧ`gRD	Q�A�i}�Z"�^�B���0M��]�.�z�6���B�I�4����hǹ<�pL	s�I�}�B�	&��ZO��f�K!�E�"O�E��m��%3��æǉ�V�x�{u"OZ4kCh1괭9�S�/��Q�"O� FU �(D�g�����*	�v�z�AA"O,�	�3+!L��!JC����#"O\��7��!��{s�H�Aט9�r"O�)a��kp�	�"�*��X�"O�|�r��g��RUbp��#"O�K�'-v�r.��J�h!�"O�p	/�����Qzd��V"O���g㈂Y�
���a�5Q�� �"O�q�7Kǐ*���E�\�_�`�*e"O�}	 aڝN�*$a3AM�w�����"O��"�1t`�4�76�b��"O^�Ń
$'���56��!�"O�ܱ�j�)X�pڂO�	�>�§"O�(�I��p���틫P�@�`�"O��6J z��XT&Q�I��Y�"O�Ց�Z# ��U�Q�@��2�"O�0�ɏ6m���ԍZ�׬��"O�(b����'o�G$�$�$"O�`;0�%�$��Y�2����"O����W�Z[���$�@�P��"OJ�3r��e�&�#E�![�@�B�"O6ɚ��J�G�Iye�
P�P��A"O��I�o�5����3��F���X"O� �L"4�p$\#K��q)�"O��� �S���g�V/G|Q"O������B��9�B"J�_�����"O|��gM�akVف$�T�m�����"O������m��m`���;�,&"O.���G4(_؝����O���1�"Od��bF��z<�Za��tH�5�Py���-�萪b燆���:�L�H�<Q�-�);2�>�6,��H�D�<	5��	�@�1��hO�t�D\z�<���%k���q���iD� 2��w�<A��� L
@��cm٥9�}��cz�<A3�D=z�e�4���&i v�<�fΫ ��e���	�T���85es�<���L���q1N�8m�!3���V�<1�C�7S)X	����d��<���K�<I4��ڐ����
���MථE�<Y�O�?F#P�0E�Ø2�A��@�<q��M<,����t���t$�d�<Y�I�"ylu�E�:��d�2�VK�<!cnC/~+��:c(ԗ/{�}��WL�<)���lR�DKU"J��Y���W]�<�k�7Z��a�HJ3x�$`�<Y�.T&�c�Г<��0��\�<F�J	�)
G�[�t]��SQ�<�Q��/@�,��C�#�V�1rg�K�<ѦB0 ˊ�Ӑ�����I�s�<�C@'��U��F
z	�4�t��U�<����8W-��`��V����)K[�<ӆT�y���J���TW0�+b�<�bȚ�F�� F��(�Ғ��[�<1�O��<�x�oښ9"m���-D������  Z�5��[+����� &D�$cPf�?7�Ū�ۢa�ڽ��i#D��3dR5/J� ����4$�m�E#D��� ��o�Dl�
�-0��۱�!D��/�O�B��S,��N����q�!D�� ���P ��H�,]�=۴h=D��Y�LI!W6� ���&B�0ѩ�N:D���ǌ��fq2��#	�;m�R����7D��r���\�f�!֯C%F�y#�5D�� �MQB"�<p��\f�o�q��"O� もX�Z�V�C�=�����"O.!�A�r-jر�Cȑm�r�"Ot �
��c�y`�YlW4��u"O�@��AV�="�1`�&��)S�"O����ϑh�r��d]D�j�x�"O�Ac��i��7i�#m��A"O����H��nX�"&��(���)w"O\U������O::���鋎�!��טP�ʀ����2d�J�����#O!�$�h�h�J2�I��DXI�H�B!�۽+���A��&_�6�g��!�dB*�CS��>=�呥���a�!�B!=B!	�ғ��r#�Xx�!�ҳ8����v�^�?���bb�E.0�!�֦;�$��W��E�BA���!��S~K�ʢcD6	��=#�τ8�!�$��a�՛�⛒k�D�A�
�P�!򄁣>T�`#��V�={� j��W$	s!���C�Z\ȣ�?zF��	0C� 2b!�d�������U)`�K��W!�$�/K 0���r�p��fO!�D����D2S����\Yz���F!�$?�4�'ǽM�: 9
B��!�9?�8����e��T�H�n}!�$ҚJ^咴�Ǒ%�����>I
!�یT&��24�_�s@}�fߕ(�!�G�[��/�%�h��1H�4�!��z�Ȣ��_�6�r&���!�$�iz,{Ɍ�x��
�BO�Q�!�dUL��)�pn���	��ʼ! !�M�t|�����]}�x���(�.
�!�$эC4$ "�/�4bH�4`1�ΓB�!�HN*j�a��I*QAX���!�$�� ��	HD�[3����Y�)�!�	�H8@�H1$L-�H��C��S�!��!`�J%:AC\�PO�y�'�)a�!�䌺R�~<�&D�;bLT���ad�!�D�4`C� ���Ȫ#Ef"�AĆ�!���wOb�� ǋ]����J��)~!��q�n�괍��5�*�z�i���!�d�V��<h�ϕL�j��H�!��Gͺ�ڠ� J���KD%!�$R>]���3b��$:��*!򤄱w�
Ɋ6M��,� ��G�?>F!�l����0�N!�2(2��(!��+RƸ<�vb ��`;�gQ�&�!�Dϥ����E��$��b�gY*|�!��=��[Ï��n��vlV�!�䁦dL\�ÅR�\�\���L�u!�פ&�D9 �Ҟ1���c��1xJ!�$S25��AnK#�岓��`!��H7��FIN>q�+�L�v{!��8EM�ؠ�EC�"�j��׋�3�!�dM�8!H	�#�Q�ЪN�N�a|�|��	�>ZL\i�O2��ASUNC(�yb�ԸP��8BP&˺+��:�$ѽ�O��=�O��P���<O�>ē���'���H�'�T�:&˟ &g<1RA�� ���C@�/�S��yrŃ::@P�A�E�arֈh$/"��x��8��:Gg�:̚Y)�;��	,::a~¥ߜ*8����S� Iѥ(�ð>QH�D�b	�4w:i�6Ð 9Q6�!(0D�(��FYm:d
 E�0� u�#.D�� �T
w�Qb����k�%=��p��"O�x`���~(����&mlb4�8OD➴ç>��i��kD�=�u� �ȩ�ȓXp�Lͥg��	�ڰ,;΍�ȓ56�}2���O(Ta�@���|�|T��$�d
֮F�@E�H��i�|-���p\[��&v^�x�P@�C�I
9x� ��Q�X����<	\2C�	�U1 ��Lg\�@��/��7� C�	�^���S%%�7~�rWI��s�B�f}4b�G��ySMD)B��B䉶i*����8m78�E� �^B�In�8��R����,��~�&B䉙<��Q�WI�)��9;��B�	�i<T���N(��hӂDՆ����>��'�.�aը�,H���[6�U0��d��'8˥NP1N@��!�?y��Ũ���8�':�\)��g�,)�ZhK�Y�M
Jф�W�%�P�	>_$�T�/�|��x;֔���5l	"q	�ؒJ�ćȓ~�$Q4�Tn�y��M�#g#�a��&�����&�T�q��P���ȓZK ����6�J�"!'ɪu�0�')�}.�*���ۃ�M�T0T5��@6�y�#ǝSf�hu��J�"�:�j\�yQ�hM�S&�=�U�5 Y��ybߨJ��8i�� �H�T�O0�y���S�r�a'��7�а�'�/�y2jJk]��'h"��@�E�ʐxRŚ�H[�q2M��<ucT�S +�B�	�M������6	S �Ū  �B�	�B�	дG��(����-v�PB�	�@�v!�0G.�������S�^B�	�7��8`�/)�4C���@m�O����Ǝo�pUV$V�d�YC��B��O��􄏃^�$)8J���d�:��/�O��j�&P��T�:�d7D�|;����n��L��T�t��t�F�3�G���*§Bh�y���N�"lR�ޣRz���EV�pAVM&���関 �pO�A��L'Q�"~���G/Q���f��$4"�T
dIÞ�y2 � j�Dp���1��;�	P��OJ#?a�'u^��6cV't�R0 �j�)�nD��O���$T�]ތaR�!O>@'���F�+mm���'&��F����((P��!��*�И�F�Ǖ�0=َ��}��D)�C�*f<p�V%$��B	�?�
�Y��2RC���d)+$.q�,�%�|Gx2� .qZ�
�.�bջ`&V�t>�B�I)#rT����(WD!B���4h���O��=�}�3*�4p`a:�a��;�d�2��O�<9��Ҟt(2`�!��#	s�%(@�V�<��O?�����HޢG����3\G�<�s�^&Ox��*�B�¥*�w�<q���b���� $;�P���Tk�'Z��h���*�'�u�4�kԏ�I����G�a�'��x¦��b�R`y�L�e�����D���OL"*5��x9d�R �֗'����֎�զ͗'��|b�,?��8KQR���R�!�6�ē�p>�2�H����,��Qd����n�tH<A���D���5���CrZ��w�I�x��(O��=��k�ap�Y�r��'���Y���`�<�@͌�|�x4(���d,�9�2aTW~��)�'*��:E�|H�Ex�^�T.Ez��|2QnM�'3�p�댵}�$=YR(;D�� �#s�͚~M:�(1�:��y�"O��X��܋'Wp)�f_�-�,��"O;�C�&&1bd�B-$��0%�PRH<y$��&/B�eY�$�r��FQz����>�l!K2P��G�.g����^y�<g@Q�@�s�R�u�$���v�<a�D�:c�,$څ�L�6ج����|8�X&�d�FL�}Q0�\7k�N9I��P�hO?�d�O���S�O%�z	HWJD�-xQ�dE{*��uQ6jϺT���,�$J���;e�O$��$[�S�F)E���	�����D�i�1Od�=�|��"�4������  x�X��C�v�<�5M����zb����B�`WLyr�'a|R%��T��Ȑ1$�6x<k�%@���D+�OrH�&J�A�X�OW�*��<"��'&�O:Eh�@���������*'%@xHp"O��[R�)�0h�"Oȃa�	JOڰ񅢗�)��� F"OV<�n�e�� Î�i�(�p5"O>Q��/R&�� �d�L� ���{�"O��'�|��c�I�)w�D��"O�,�"�[�yC�ᩀj�?!�  "O^�B� �}����� %r� }cS"ON�R��$T
����aW $��<�R��G{��Iܺ&��pH��U�T�;,�0i~!�D��������3,r���k�^2"�O�,���R�Ҭ���܋�����"O��KE�Yhfa{�F�'����"O��
�1,X��
K��u�"O��kUj�M�9�̤<��`S'�'Q��u��� %c���-<�<�Y%L2D��S�f	@�L��oިh%zi;�0�d�<�~"�i�j�|z��%S� V�S_��zC�ɮ[� T��P,����U�܉��{5��q!�~�8 �{��I�>	��GJX5�Ə�.8��t+7�JS�<�!Rk�d�[Q̗'=H�lWgy��d"��?�{'��%`@��珐i	���q�.D��{Q�ҍM[��#�O8V���.D��BB�2LW|�l	<{�hI��,�O��ɇs�0%����(<le���NC�I0q�5a�ċ.;8�b�B�w@�ʓ�0?q$��>~e8����]�x�
iӐ\������O�[V���(V�9���K �
IU"OVm��e#�	 ����b �l�<�C	�$NJz��n�+vҾ`B������xb�^;n�l�s!\�5�u�T�X!�y�j�8�:���)
�H9#��y�(��	�عцͲC,�y9򭐒�y��!<1���fgD@�̈!oV��yҫR�{�j�s�d78 �hQ盬�yrB�W��fC=�����y�L�D��}KŤ�5�S%���y�ɇw���Ce��&%V*l ����yR+T8{L���">��o
��y.�O�
(�J�9m����F ��yrM�-׎m;e�{%d�a���y��Ӌ��aui�������Ȇȓ'������_�V�1+A��n�z`�ȓ7���"�݀1{`�ܖ 0��ȓxKx�x�ȗN]>I�Pk�9`,��ȓ=�|ԹuB I�n��0�U�D�ĉ��S˚!����[/=�b���q�����]|�ɅEιQ�B)���怅�'z��3ȅ���� A�-�ܨ��S�? �PRq��3����b���}�"O~|��ʔ{؝A K��wDЪ�"O	��eS1(D4�jA)�&���+%"Ofac�`��A�3/\�T��!�"OJh�g��H�09hBM�G�hErG"O���d%P�9��wiޛM��Ńg"OXؚPE�)h�&�AUg$=�d�I�"O脪)ħ A�]�ц^����"O�x�W�Ƽz�}�#�P#.t�$;�"OP�;�F�9^�8���:\q��W"O"q3EGW��(X��L�/ώ�bA"Ox����:��:�d�1V�Qa&"O�4�QIK�M�	�X�Z_ɺ6"O�\{a*@�t.h�@"�1H�5��"OD�j�Ǌ(6�D�ZWp)�!"O���πI*Tu�#�@	(O�tK�"O�=(�"?,���XG���8=�Q��"OL�y�5L"��
!.�,g�^y;�"O� ��Œ�kZ�8[�-A�_zj��"Ov��g�W%S(�@����j�@�V"O���͆]|�؀�A�N�i�"O
1�tJ^`qz0;!D]*D�T+"ObMDo\fZ�����@&��&"O�y�B	��l�Nu�e��=2��HQ�"O�X�#^,���� �C�� �"O��5lN�,�����D"O ��D�<|#����䠲"O�,  ^�! Հ�/2$� �"O��V` �]Q��2�\c�"���f
,��eQ/��YH6�'��=Kd�B6C #ˆ�hAK�'JP]��������x?p�	�'D؜X'g^ <�(��[�wy��I�'i��k��ެX��lP�O�_|��'R�5��ÒP���#*׍z���j�'���{�
{���c0�
j?D}��'���j7�Ӈ:pʘ[���f-�h�'��qJ���E��!.pP| �'vl��B�\''.h�)QF�'& �y��' pX{lN?�a&Eƴ.���	
�'���S��S��!�U�/O�c�'-��m4�����lЇ'`�Y��'������DX�E�!'�� �+�'�����iʇY\���a��O�����'����,�
�::��RV̰}B�'1�Ek�̒�N(IÉO�Mb~��'�VѪ0h�D�h](b�A!�x��'-"m���G)許�1d��"&萐�'bbűG���i^��`��MZŊ
�'\���Rψ]+�,� њ_^�)B
�' (�p��l%��[0��
` |M	�'6t� F�F/�~0�w.�jH4���'%�A��K@�9��o��Љ
�'�T(��i.f|� �a^�g��, 
�'��Ӗ ں
3�T	Tj���	�'�Z�QF��:<�
s�5W���1�'��c��rZ�%�d��^(:Ź�'� {f+���U��%X�b��
�'9\%!����.�fQ�M�,'~5��'(�,0��'�X�K�E�
6Ĭ��	�'-����

2�N�ʴGۀy1��	�'d�x�s�6N� 5���A�N�pQ��'��h�h�P�v4�C�B&���	�'~j�`f��?˖y�s2E�ƍ"	�'����CC\	S�FIw������ �	�lW���H���~���ȥ"O����ᚺ8�`��"�",r�\� "Ot�JY�\�����ͅP`
���"O�Y`���28ɰ���3g��H"Oh�#'���cה��F��:��,�"O\HAmХrvy�ߺM�^<A�"OĄcg�5c��[2����Ve�<ɖ+�E@�(ҕ��b��;TM~�<A�E4ͶT�F��o���O�a�<��C� �X����0�U��q�<IkG=,��t�^A�9S�&	Z�<A2���]簕{�G�;��r2
�B�<I׋ݳ�+�7*� Cc��C�!��Gb�YjC)H%XU �ɄIy�!�d�xФd�7'^�uxx�4h�5k�!򴔔����ky4�  �	�Ф0�'Y�F땯UW"�@4�)��'���{��M~�H��	"ʘX
�'�4E�f3!��@!�kړ��
�'3,��H�p(�}"','-�9��'��	IfJIm���{gbA&L8��'�t�8F��3*��̢�I�'9$y��'����
�:Ocx�� �4�'O��B4�<E+��mWF=b�'P�d���H�qs ������U�J�4H���/qO�`�Q)l�Xa��؞l�,��U"O�= �I�Wz�k��;L���"O�\�Ĕ3��9bC�s��3�"Ov�W�.p���:F���!�>9z cG�q$��&Ä����!�)擐	p10.8�R��W��#���p,ƭ0!�.�	���O�`��҂
D:�y���G%ov�I�nƏ+,�J��4R���x"�R[�:l���ͅ�f�T��O4s��Ŧ]� #���o�'�(m�UD�o���7���IS!��QF�Ʃ�=|q�4F}`}��5� n]
��p ��;ղ�p1h�3wlP:�e�
��d �,�h�v�0dg�:5,�Χ"u
�y/�*�L�c��Q�I��?!#�O�I�o��/�@�sM~�ժ�<��m����{��	WDړX�x������%��hsC�)���'�')kd���U�j �"�bO�X�6M�@���!-�\�J�!1;O?��W.<�pukJ�b�
��¡ 6�I�bS�V���!�� �/�  S���}��}�^1*b-X�L����FN8�M�r���s;�����<�(�;Gn;"�D��uO;z��s�Ӆw�s�H��X�����OН�.�1M�:&J�*Yj�qŮ�x��5�@��b�����|��.`����S�4���X�N��'��1 �06��{�&L� ��6>n���� G0#��O\fY(n� r��Q� �s2���'��(!�s�K��ߒ-VryRn��p��y���r3� C{܍ �f^�5n�ɨ��3d��7�|����g՚ӧ�T�gא=C7�P�>����r�S�����<�&h)�n-[h��A��� -��T���Oar�0��ܬ|~�� c�ix����c��	 ����*�2C	���5�N�}�Ė�T��%"ش`���pVc��b���X/(S�PL`9�8Qi���?y�ٱz'T��,rU��+I)x�*1�E�[��` �V�Z�����g-^��FfB �2ȢE$վd��%@���m��3�a	5@Ūlz�hD2d��]ʍ��D�'�
���5�ӉRQ�	�0OT>�2�y@�4$�Dޱ	�TͰC��d��	�s�Bo|�l��V��0��(�O�z0�#\";� 쩔N��V,E��O�I�si����u���rDJhѴ)��F��B� �2^��m�R��k� ѳ C+ `1�K[�-�,Ո��A8 &�R*���~`�c�Ĉ0�AC�@|����� dʓ�ʯ0Bd,��%4*�d��'V�Ɏ6 #�*2M��b�(͛z�Z5	p)D6�V	���!5�ڰ��' ��i�`�٦(	�`	~���#����To�u�⠀
P���O�ͲLT��2�be�ׇ�5�l]k� S��,j8���a�C�k/���I�<��C�7�I�q6�8i$���qp!�K�B7�%�Na��i Dĩ��/R���� �x��a��9j�SX�0���S�K�P!�P�X,%��Y�O���1�M�w)6}���1�l1i���J����"�r>���ɬ$�(a;fɕ�X*Z�1���O�VB/H݄MZM~�=q��I>@jd��S��c)��1�@����V���g�I�d���[�?���	�|虻&���⁑�:Q�9C��L  �\�i1(�<"��#�߳��=)��ܞtVRQP��~�-P"9���)�eԔ��4m��<YtG�~
p팓�x�$�<!7��
�ب���!��0t�xX��%��'r>���%�&2�l��A��*Ű&��=U�PB�΋7>�pえL��|J,�� �T�B'H�| Yo�%2��0����@��%��e���ǔ���	XפȊck��{�ԁ0ʆ�yZ�B�	�j �ŒVI�`hX*� �OblHD.��/�4!�F�9}J~���̹x-<�j�EЄ�Dݨ��$K*ʘ���#|OhD���aYxi��,�5�����b�2*�eW�F�O�m0L~�#3}��ƛ`j� dEĕ%�% ��J��U�7��"~�R��1�J�i�� -��t�æ�*c&�;)��:�Ea�;(�����P�r����s5<����y2W�<1G�|ʟlp��#MX}���WO8}���1ڄ�"٘'	�?��|���'��WԲn���QG��9�v4Di}��zX�p*�Mǌ]�dH[���R�A��'R�v�Ѝ{��O;f�d�R?A!W��c3�^�DӾx��M�^ �#�'���'m����`�I�'�D�[)@%!W%\��~�X�����O�8?%?�!	�a(¬���Y�����Zf�ɛP�X%����P�\��O�@��b��$���Օ,��Q�0�Oƈ�觭���g8���>LL^(�"P�K�(x����X�!�v� �=�O"��h"ЏJB�H�dm^�m� Hx bȈ! ��4�t�iݱ�S��83�!�~�M8#N�V�`����"D����F.N���0I�5V����έ>q%%�O8IZ"�Ռ'��T"rD]~�(��'��ϓF�z�����+}-��P�LԳE �ȓq�:%�GmS,q�` 2C'�1��mF|"g�O����*��L�H �cIS�h	�'Nxq��`��E��A2"F+�E���(��<E�eM,7*��s�P�mL��020!�D�~C�����4v�.�����2��./��}b�C�[�HT�A�T�:T���	�p>Y#&?	2��7/tj��wA��3�|(�b�9 ��y�R�6�y��~���vb1pAcܦ*1B�X�-�>�O�Aڏ�?���C@<N{D�X�%Y)�))�<?�Y^�|�_�-4瑴�i��E6}�l -��K}2�� ő�5KIk�m�,u��9�	>d�}S�D0�O�<�P��$kt|B�ΞvX�c�i�p��ɻ{7�e�箍��?iҡ�w�>0r�
���E�D��P�'($m��FOb]ɏ�4H �C��!� �\�wf�����q�<� ��(5��`� 	�06j�r2f�P}�'�G��H�H����`C
y���U�`�PS"OrD�G
��I،��C���Q1�O�E��&ԯ%����9xF��b�^�IA�DZHH�a|�gңBG�T�%�\<#�r���Ó'{��H�8!dqI�{b�ќ�� ��I-WKʜ85��RbrĒ�ƌ;?�㟜a� �5Y���	!*ZB�'Z�����jZU��� ���.HTm�nRV]���'�LM�qj&\.t�A@�S���	Ԗ��H�e�G����p����W�3N�O��PQ��.:Ѯ��	.kRd�`
^x�<���^��<Pkժ+M&B ����1���R��Ҵ�� h�l�B�)���)�C���h,K�|5SY��{�i�2@��%��n�A�z,� Y�%��`שU�7����GR��*_e�A�-;��$� :�kgj%r���M�2=�O��agN�x�)��4��9~d��P'"����go=�Q�$��o�a�	��6�0����. )Ұ!T&�7l;�JS����B�[yb�O�0p`g�I�1k��OHa� �+.�iۂ)�a�0P��,D�9� % ��m��V�N5����O�Y*�Av���T���	1.�:�:ӡ�i��Z5`iSw��\S��{��l��*F�[f��k�|Ԛ�C��wG,(��K���\@��-���z F�2`@Lb�3Xz(PRqM
+�L<9���:¢<�`�Yx,XZ��4`��I�a��芋g�Z�[�@`��d8��B�9x"V��e͍� �2q˔�p<Q�"56�b�� )'2Cly��ș3qxxpP -D���PbôoX]�G��_����E++D�<	��S��tC�֜2��I���%D�\&lϒS��Z�m�-�����>D���Æת#+��Q�-˯&/`i*a�?D�D �K�����Vኄ|:���/D�X�׾lQV�k���%1��!��,D�� ,�`�gC��bdB�8
��G"Op�[���C�4l���`R���"O�����-}ȍXuN��A���"O����g�- S�\�Ƅʮ i�*�"O|X�F
�bZ��z�CK�b���E"O���X�E!�Ѩ��d��I�P"O"$ Wj�k�,5 ��?����0"Or��Te 5@��.��4�H���"O�ٚ5���~G6 ����h��bc"OЍbe�H�{�.���c��:�"O�@��]��A�e�4m,i@T"OB��c!gQ, A nN�[�x��"O��*����T��c���:@�^)(""O�� ��Y$}e8����a�fa�"O�I���˔M
�� �Β�u�j "OtM�3%'�(MQ��Q�ul�u�"O�����xܫ�k�Cv�b�"OXАB"��|���jDE�a:�"O@���lй1g.1`��&;"�� "O�)��J�6T�)��364N*�"O�P�G(�7w�ܘ;��)^U��"O�Ѣ��'�d8�p��?d<�w"OZ@irJX{0E`��@C��:"O֠E!2~wj�("��yG �B"O�t0� P�54"��v�Z�M=���"O��k\�$	*r���"Xf��"O�$��eY?P� �	1V�""O�����5n`ڢi��PuSq"O@���F��Ըb�Z�R����"O&E�ч�8~���Q-�$v|�b "O���O/:�����-� ,�S"O4��b.��]Y��S�`2p�qi�"O&�+!#��II�5��抪i@���"O���mG�	[��O�0Z���"O2l�#�HU�^ypG���&��3a"O�y[c���8�d� #��eW�t�t"O.��-D�Bd`0CL����V"OD�K��N:#'Mу�W8ؤmq�"O\��E揁˔�C��d�<�Qg"OڼJ6U L�	�i�?� ��"O�m�A��?u:�����F*S��0�"Ob��0� �S%lir�u�&DQ�"O E�k\#OM��LD�J�ĐH�"O����T:C�tͫ}����"O4�#�µ�l@�B�řz�D�c"O����,NcȐ��j�?�䈊�"O��1Q�r���Z�cNO4"@�E"OJ�)R�"$J��EaF$��"O�h��`ش84E� �˦m�X"O&4Pv���/JY�e��b�\@�"OH� ��Ǝ<��Z�̦w-`�ap"O0�� ��F�9ᅋ1 ��"O�-2�H�_��H� �
�>�5`""O^��t)����ɥ句i� �X�"O<��Pi�"��$�Τ3�Uu"O�|1B\_������iJy�4"O|h��ƻD@�]+�� e�p"Oth��(O�n���HaW�xĶ��c"O���� �0�&(h�OV�R���
R"O@B�!L&�i�娘�`���a�"O�x�A�
%��Ѱ/h5>q3$"OZ�5�F��9Y7��R5���"O��xUH7�(��Oɹf?h�"O�(�2gЛz�i�0mK�L'j�cQ"O� 
�0���O"���&j��K���R"OHj���"��ժf@Zpa�"O�͸3)�<qo%�c��A�̒
�'M�ab��U�1��XR+ڵ�0X�'i�H�d��K�d]qAJ ;��c�'�	���Ee����,�:�1�'�n9 �	�*n�i�� �^l�
�'�
��4��!ے�ZT�$C
�'����IUc�کirJ�L�>9H�'�����k0�6�q��Ep^i��'ɴ���$4�≛�N�sJ�B�"O�xx�ϒ�����bm6ogܡ�"ON)$dǇ$�B�q����|] �@�"O��+QD��J=��uGՏg`t��"O����[�x��l0C�1!!��"O. �t�PHm����B$̩�"O�=�!�T#^F���C�t���"O�Px��ɛl���0�����p"OBT ,�P6�r`��(���a"O���ց�$o�J�LX6zeP�F"Oz@���6X���넵
_�y��"O��r��_O��(����$9NQ�c"O���E�������w� �c"O�u�3��M�I̚̄+"O��Z톇wTTB��A<�A�"O����EZ�^U��zȷXf�Yː"O�mHB�M��f���1)E���"O8����ѧ<�� ��.6 ExuRR"OR�Z�c�
qH�ieM�"~a["O��蔆9fy����Y?D���"O(�;ą�>%��U��+��p�"ON�s��
� ��jK�8-�P��"Ol���"`*��!��zJt���"O�]��F�NԖ�y�,?`� ���(��&�qO>�S�L� !�LH���¯j.���1D����n�4+ex"D�U"8��:�d_P(,��$:O8�"�C&ena`fm�.`��{�'ndeb5&�^wd�h�m[!�Q�$^�)�0�%�J��`�!�\%6� �0vj��3�9+�c2�P�&��a��P�@����8�'�9����p���)ZRmb"O�e8"�@2ƴ���F@���(��Q�p֥ǝ0��(�>E����s���zÎ���E�U�t�txׄ�&}���"~�	�v'��sAl�&�<��������ئO@mJ��� S#)%>c� �JC�e����bУ E�|#�{�@H�
�I/9��	�m��Ъ�	�4����H��:��	�U�LT��C�=��aI���f�~b�	S��ιq5�d��9��q� B� �.��D��I!o$�S�`ѳ�Oj� ,�u���IQnX2��q�'���y�O��e!�+Kb~�0R,9}bF�|���M�d�Bq儹2��A��FUm}�Ջ.+ԥ���
V�ԟΝɅ�J5�dU�c��&����$��+��	vHɠy_�|[2oL�d��J�l��峟X�u�O�Bk�][2�ؑ-�x���$E�$� S���G���Й�h�iI��F�;J��
q&�� ��s/�����Z*'���ɋc�`�QW�9�0<1���K�r1/�<�  ��
��*m�W١��К��1yצH��� ��V?I�r�F�L��@&�i�
�:v�����05-n�XZ���X-ts�3C�4� `6r\��K.T�>Yb��-K��d�4Y�|�"lR&`Ւ0$�e>zX�M�ȊEQ?u:S#�&u4"U{��ӡ�����=?��n�Bh����  ��(�So\�5?�b��2�|aA@�J��T�1CZ�u���`J���ɴQ�Q>��(#N�c.��a2P�,�4�����G�TL>�@g�'/�����y��d@��I� ?�s�5O�`f�@�i����6n�Q���o@"5�5Ǐxf$t���4��Vds?9���,V>`�͓0��I�d��)/.:	G�DZ65�ȓ[�܄��D��}UF���91>lڛQ�����ʩrU� �1�'�����J�X��$x����)��sד=�t���
:�p�Ǧ�H`�D�B'W�Z!|���J�z-�C�	64Y�#dߋ $���b��?v��tsQ�F>ɠ)8��3� ����̎27[d�ң�W#L5��"O�Y��ޖ ź���*H�?*:�AF�&gs�q!r�>A�l>�gy�h�����$�߁^r���hߊ�y�N�#�N�aPm�?�P�P\1aO� �o� ߸U��|� �Cƪ$�F��e)(_:����.Sdhi���VE��$G�9�H����/0c@��+̓}�!�F�H]4SV�S%�du(�jѸ?YqO>�`5(]�)<�U���I��wQ =��H"�	J�j@�B8!�!PY�=�ѡA3M��-���7�|:奟��dm��|�'�
P����/('�]��
�ܠ(�'�%��[�D1��Z8����42��i%���p>A�60li:EA�G�F�pg�R��8`�*DVq�	�$V��iV�L2	������.^>|B�I7g!P���T�(~ ���ܹ"�PB�	�&n�mʥ�ԫ*t��A.;O�B�ք�bǞ�v=$1��.v��B��B�Hx�M�}+�\�/��k�<C䉄m� |�@�M\���Q#Q"v�C�32��آA���f�l������B�ɇhNʔ)���Z�l�4N�C䉷D$�X�ᎆ(�։[�Bd�C�I�a�\��!�]Pt��f2ZG(B�ɴ<�|8�/V�?Vp� j-o�VB�%$�z�:�"��E��sjзl�B�I1Q�~����	�%��m[�dЏ(�C�#hP �$G�@�2��O�|�:C�I�J
~=����f����).O��B�I#�@�RAR�w�����V��B�I<f���ᓛy���D93K�B�	�A��������P�co�'��B�<>�������6ᦈ�r��rp�C�	�1�F@cAH���̫@@�;lE�C�	�B����dǝ)L��T��k�bB�I"��hR�� �����cV$;�RB��G�Vxz�oTEz
eB1���sl B�	�(LPM#�Ʌ�<p$&N�+�.B�	.\I��v~��Gӯ__�C�����&��.)3R��cB�j6C�	���H����p���E<+HC��0Gi ��$@�x̂�eU�h[�B䉇(.(ik6B� uF��w�[<�B�	�G2P0��?m�\�EN=Y���!4���x�l؞�PUhV&1�H��Ȓ.y�I��0�Ov����l�"4k�$Zt��"�ώ$��Ҁ�=ZqOZaP����0<	)Ž�p%Yb��@��B�S��pA�Zb�x���B��LRy���h�4SP��ׄ0`�6�xal��G��b�N�@��-�������5���^�x� K�d�<y�'@��5����ӧ��,�t��$��]¤"���y�nTG,�-�'B��X��GBZ3�?a�bY�x*��؁���s ��'�\XqC�9[���+��xP�4X"쳥���_�V��d��XP򔚥�T���ytQ�]�bՊ"�V<���ap�ל���-����[n�3��&�q�Ѐ��<��pX�eN�o�t�ā�M��K�5���w�.O�5�Hӭ><xh���	�<h7��x� ���':��y�D��7n���0쏱O�Ĥ3��bF��)c抬���%iFf��.�8�K�<K��T,���C64d��rb�b�<14j��E0�Y���&=���[C�[ݟ\IT��}0\��λ7&��@��Gџ��iX�&�h!s�P�rաb&Ӌn@a|ZIP�pR��ȱ-L`�S+��[�VD�BL!w������&��ɘC�bu�g�N�3�I�S�Z�p�k��[ �#�F�[$�<�R�^�x����=�b8Kh@2>��l�&c� �5렉��5���ɐ#�\���e��d��Nƻ�p<y�N�BF�c�X1�Ku,�ېΝ�a(�m��;D�,�UD�j&N��"�[u�e��:D�x�Ek^�sk8A#�)�����3t�;D�� R�q��;;�x@0�E:�()3�"O(�@���<;X���C⛭�*�!�"O�tٖFX?���(�fl ��"Oz�B�.�$z�:(�R,M:vg�|C"OZM9�+Ǽ}�Л���fl�MH$"O�1v��:>(Ř���Z�Uja"O�������|��`�"��XP@��A"OҤ��n��D|h�i�"BS�x�7"O֜a���H�a�!HtX�"Ot�"mݝ|��*'�!$r�`f"O �(ׯ�m��l��a��`-���v"O  �7�މf���q��!�Mʕ"Oxe�סd"��z�LMy�t�"O��2�5>q�I��j1�94"ON-�G%�|�X��Ag�%����"OR���aǻ&���ӷ��'2�A"O�t��'&�]�h��S��(	�'��DY�,ȭu!d]s�E>V�x)�'�
�{�b�{�������Hz��J�'Ь�ѧ�A�O[(�:�JK�F�"Q)
�'��$$���i��u�T� 	i�@�	�'���(O�  �aa�
�`��	�'E��
�ٵP���0�h�X��	�'��H�E���/��`)�N�j&`�
�'b}�s��2b��+��&X�l�9
�'$s���K`�@2N[�%�nD�	�'w��(�ND?ؐ�	R����	�'�y�r��%
ma�N� HX	�'���r�Ι�K�q�孎��`�S	�'�$,�f��3(ʙS������	�'2��K �=Ft��%�		�'}�j2�^"}Pr=�A�?��y��'T6�#��U�HF ��aJF#	'4���'������-\���!��Pu�8z�'��yt ��>�Hx�"�Z��[�'i.�8�fD�`l2d�"�̐R² 9
�'>ԽRa�R ��aN�A� ����nĘq��1�a�L��r�%^l�Vm�%��a�`|�ȓ/�A�b*�މI�ɡ3�����OZh�p*_�z"h���3I�ц�+�v�8��Y�E�L��T�/@<�ȓTƨ��B	OX�뢋� eTr��ȓB��-%�R�H� ��-Ah�����_H�1����
c��:��2h&݇Ɠ�>�����7OL����aN��"	��DN9� �͓�Z�xx�Ԥ�)䐧Oh�i¦3qؔ,��#� ��8R!�V&m�5�m)�)�T�`P���H��=Rê'>bJe�A��O�?a�B��Ej��J���v���^r�'*�#=�O��y�` S�m_��0�$����{�")\O�Q��`� ��XR�D�1����"Ol��ʃ/*�#I�2���"O(����)v�
�	�+N�GkyB���@�O��%C�葱h4:�����%���p���<9��I7K	Fٳ�Q9dIzt��ŗ���"S�Z )� ��r��<!���y�j�]�����+#.ܥ��'t��l�D��l�!�dVX.�q�[Q�L�S,��!򤇭K��Q��#&��I&�<'g!�D^���Y{1�1s+d���K& !�;=� ��E���M��'�@�!�-[���)֦�*��h�@���!���**�X��eA�8>�PTgןr�!�Dӑ�$8�.� ����GA_(!�D'���cGBɓ�2A��z!�D�`����	Ql���Ă+8!�� h̚�X1@; �h�oO4/&lqj�"O�h���5�z=rH�M����"Oz܊"+T���!c���JR4"O�d���K�g!�mڰ���| �h�"O\����5+��Ѥ@�t!
�"OhP���̝k������"}Ėl�"OVU��^��D�`�
�"TARu"O*\i�Rl���"���X "O���BǶttq�h�N d)��"Ob��tm�.J@!�։�[LZ�)P"O^P:���hU�0��֒y!�qT"O�8җ�K8����-�?/l�L�7"O��u��2�qr��6�d�e"O���S�ց���Ǡ��mz�"O�C��u��i�$��LH��W"O�(ţK*�b̘�IY"g3>�H�"O�����;׈Q"c�X @#�u�F"O��,�L����C6$j��"ORDk��P(^�~�8� ��,"Od$2�$U%h��qt�S �9Q�"O��L�3i���06L�P�X�"OF� ��2L`IP�B�l���r�"ON(A$IM�(%* �%V�
|��"O̳W� ��1�9�pd�"O�K2	��(��T�$'Z+~����v"Oļ��&�Jp0�(R ]��0�"�"O֔.K0ib�@j�l���[�"O��ff Y(ڠ ��R2l4���$"OڽȂ��d�E 
3d.��C�"O�QҨ�A�dYg�0O$����"O�S����|"�J,YR�J"Ot31�Z�Eh�X&'�3*rip7"OtQBv�@�\RDC9.�ݢ�"O����@*<�`��!R,<e���"O�m�wU��8�8��R�Wyh��U"O�i�R��*1`mp��Ʌ
��A""OДab�]��E���G�R%��A"O<�1���@��Ѕ�3�l�"Or�h���.̰Cfo_�h���7"O� ��@P�:���ֈ��e�8Y��"O�m�b� ��PRE��C�4xw"O~	@�A�~�8 �]�/,IYD"Ot��j	�d��Pw��ǘ�I�"Ov��Ck�0��9��!H��\�$"O(A��9f6 ����_:�X���"O�a �n#2p�ݑ��I�X�"O<̲��@�$:m��[3V��e�"O�Q�C��M����e�<��(��"O�I���	>Dr=�Ue
!c�h�w"O�}s"F߮p8v��,P ��"Ot�Y���*(�C#��P2l�S�"O|c�Lۊ���d�$˦�ʴ"OT�w�ܥM�N���
S Y_%��"O��Ш!tkdyGG�#E���r"O$�F�/CE�4@0
-�>0��"O��c��� 5��y���7��x�"O�����J�q�R�N>gra"O��SED	-J�`z�	�R`Z1H""O�$�sd�.{@(1*H4S�-X�"O�u��M� ���ƈ/;M,�K�"O&E��S	;?��(�L�D�f"O840eGL7QGh�r&�8�ޔKR"O���+Uw���i1�� ogX�Ae"O2�K�����f�E�I�Ie"O� ����_�n�ب@��J�v+ ��"O�����ejЊ̘�-JIz�"Of �E���rj�$�a�OrA�H�"O̼�-ԽZ}X��%�� 
2�a""O�Y��8ef�sF뛬`���C"O^����N>-�*-���A%�)��"O�R�&Pi[~)�2肼Z��+�"O�ri�g�@�BcfP"	���
�"O�����	Wi6�@�J#��-�D"O��y��G#GF�r� t7j,*%"O�y�B%C�#䁮;<$�"ORi ���*F)5f�_qS\��r����IHPV[Q �V9Ѕȓ!�5˷��,PѠ���@11re����rĩ�3�:����G�g[.t�ȓGz&���[-��tҵ��_���ȓ������	(,|�h�4xx���ȓ�N][ǎD;��}q�Çu�F��d�0�Qa
$^�"!ރ.����{�"�	�&&�2ј�N�68B>}�ȓ1T�8�3ʔ�&���$Iǚ;��A�ȓA����j��Zn���eE�j��,��>���	�H~X��a�P�C���ȓN.*���m��/��`�@B���0	�ȓJ9�h`�����IFnHL8��ȓhH��P���� ��'��(��#TT��׼:2e0.
7�V���5�ݨ�EE
>��{0@��ه�of��a	�9�nq bC�KFi��*���++vF`�`M$R���ȓ���"5�]���\�ee`Ԇȓr��`&"	��T���g��|�ȓ~���ҪQ���Ժ���z)���ȓx�tEѤ�6hD\�SoG�9#6���UҀ�S��,��5`�=_���ȓ����ĺWr FJ�j��̅ȓ{b@��F��"J��Ac�Č�x���M~Tɣ�iM` 
��p�l�ȓ��9FAS�n�lei�kY�<[4x��o�F�����V�^!��1h{܍��Qp��Pc�νt�*�Qp���~�N��ȓK�Ri*GJK�[,�K`%֭)����M��A�Rϋ��Z�ð �&����JʅY���&:��Z���-X����#�bHr����q4JΗ`��ȓ�x���	��}HC�E�q��|�ȓ.1N)�o \��`g�;c-��ȓW�t�1 5Ԗ�j#�ø mA��Y�СE�@Z(�*@P�g\܅�;�Y�����?���[*f�~(�ȓ!�}*W�V88�u,F��"��@��:���5���)� �,u�f��ȓ9�Ƙ �̿^�r�GC%hAV���_��H怘)���H�&�^�x �ȓu��	a��ƟH�"
pfI3����_�f0�d ��N�Z\)���-X6L���~���冐�"a��åe,H��v��4^G h)�R�~a��ȓ CB��Ï[�47b,����Zw�نȓSHN���kպ	��!A���h�lD�ȓ2��2f�� <�<ؠ"���Tp��N���� �E����Yy<��t�ձC���l�s�#���ȓ?cN!�F�
�� q%̂%�l݆�S�? �Ђ�.�Y3��CS��-�����"O�Q���M-fU�
��Q�@��0p�"OFh���O+{��1#S�܊�2�2S"O��c���eqj���j�
1�:�8@"O��蘰�����~q��"O�R��s�A�Ӈʰ̔� "O�L`��*^܄�r)�F�P\��"On R�`���,�ק ��(AI�"OF���	`e!Q��m"�@�"O��r�R�l�����R>b��܋�"OD�7�
�]s�)3��Q�5"O���!(�9�@%�5�¨|$^䘦"O���'�׶]lu����[���""O𰓴
U�HN\��	�R����F"O�m��o�U�H1����B�L�{A"O�xxg�F�4�KW�N�7��Xb�"O�`��oY'b$�;&�ȺzJ���"O��B��Y�e��r��7`_ ��1"OB4�Q��.`�$�61ZT�tg"O��14�P#>�4�2g�+,9�+�"Ob=X7�\<���f���"O~,Jd�E"Su�Թ��E�|��"O�a�S�6U�@ظǢR�$�
%0 "O*$�2W�Uf�[����@�KB"ON\����9��0q�)��F����a"O������aK�@�1���y�ּ�"OP+�gɄli�p�#�>k\�i� "O>�AXЌ27lTp�2팩�y���:��:@l�=�Ja���y�-�N�<<)Ì��
D��Z��"�y�C*p�ܥr�c�Y�b��VM_(�y�K�c1�L�E�@9N���v��0�y2F���1����0�pp����y҉K�o5x����4\+Vy��g���y�͖�b&��	ЌY�A����f(D�y H늳6�ǗCG�`�ܵ|bB�	�,�����VQ���##f�:ҞC䉭7㼥��@��v �(��D�C�ɺ5�z��E�<:��5N�0B�	�ug,�(�ތR���J&�B��B�Ɏ1���7�7�ɢ5 Ĥ	��C�=�U� d�����6�� �C�.3Τ� ��P+Q*�8!�A3d�B�	�x�9��(:a��/=�C�	t�S��n�!bqʇ�D�����8�����VzJ���\��!�\-�j hh'OHN�!!��b�!�4(�H��hI2	-��i�7&�!�dG\)F8�#�@6f������u�!�3ɨI���KǴ�`'�K�!��Pu�G��l��#���gr!��R):����=��F�oT!�iB&5�6A�/[o$]����2rY!�͂k��x����|�|����"I�!��V �Z4��E ������NG!��3]t�*ң�E��I���l,!��*n	9����X�2�bc��X!�d��F�|��	��`xe�`a��3�!�PH�M�thJ�NDV�KJ��E�!�DU:,�ؑYS�ϣP,�5�B<&�!�$V�_�LH3"�+���CW�J.KV!��Y�Y#z!C�K�X����ѣ��ya!�$�H�(������Ĥ�ГÀ�d�!��TfnZ�[�KC/�������	�!�� Bt�Rϋ�N�����& ���"O�(C��� �b�ʲ��5<U~E�"O���   ��     G  �  ?   .  2<  J  EX  Gf  !t  �  ď  ��  ��  е  ��  o�  0�  s�  ��   �  D�  ��  ��  �  y �
 � r � F% �+ &2 j8 �> �E dL �R �\ �d @k �s { 6� y� ώ ��  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf"O�Ya��=!l���Ɔ�b�V��!"O�!)��Y�fx���eE\z0	J�"O>��pg�0Z�2=�C�A�Hy�"Ob\B��;h�`��Ɇ*���S"O�h�T�ÕZ(jܫ� ��+�Ƚa""O�A���I�{"��qReM.v�\�J"O�I��cR�G�Fm+De����(�"Ov�M�{�Ҵ�U���F�T��"O� ��M�g��l�a��8{�Y*7"O�Z��іh��8`�tm�`�"O&ESS��M�,ɠ��b��b$"O,y0GD�!�<�Y#dYF��c"OV�Wc�6�:�3�	�C��:�"O�`y!�������3-�<�"O��!S��3C����ǇZ��\�C"O�V��vA����EE�@�J�yT"OtXa�Ǫ|�t�2&�ۥF<��BC"O�i�w��&dUj��+,1�4�"O���I�tͰ5���߷O�y9p"O��&�(w�̕Z���
P�C�"O1@ŏΞ
f�}KT��}�P�&"O@%����-Zw*�`C�#���"O01#�m�{�0Rda�#�"O� �	�e���Z� TX�؉B'"Ot�[��*Y�~����4[�h�1P"O��@�K�4Xպs-َbF�ģ"O�-��H�l붼�t,�0F(���!"O�����G>�`R+�0Zy�6"O�eXu럋>���i��wf�%�Q"O����d"�9c*��h>�`;�"O.T���T�`~fM����q)X�h�"O,�YD�#H��k\��t��"O�ɢ%b��/�P5P!m��hb5�%"O���0�φO�Z��k͡1���k�"O�``I�4g$�1шىK�yR�"O6|�D(
46�jf��\��A8�"O�ukg��<Pz�Aa`�#�h��"O@PQ%ƃ^R��p� �p���"O�xjd�j���a�ݾ
L�t�V"O�(Z�[�3p�����CE���r"O.��E�	Sn���
W)^?n��D"O����)�e=!쎷E+���"O����!,\�| �-Z�6xtb�"O ��.X������.��K
�!	�"O���*� �|�S��N ��irU"Ofl0��h=��@�D 5K��� �"O�<kqO�D�
�AۣFj�@2�"O�2���w��"��QL�.a��"ORp�2H��X��a�Ԇ	���A"O�u3o�A�dr�R3�Vy�!"Oؔ�sO]�:��@��z���U"O4�k�a].����E�j	�p"O�1`�	
 ��x1�F�C���XP"O�𪰇O�<�D�8��$m�p��"O����Ȃ0z�L	���K�(��	ˆ"O0���<�*��4bڥ�V<(�"O�m��OE SX�7$�f�31"O�x��R�8�k�]8�U��"O���/�4Q����TdN�lЌ�Qc"Ov���j�3����cč�Dm��"O��ۗ@^�?1�H��ի:�晀0"O8��M�T#Z�h����B0p�r�"OR|q5��*?��ATn�(Ta+�"O��zc��n��w-ݏ���v"O|��u�&�j���?$��q"O~4���7,��)q�V3h���s"OJ�r3M�i�[��V�ZY�u��"Oҍ�dD 0��ER�<hbv�A%"Ohx�  >,jȁ��"){�M{�"O�(�b�Aq�tQR����]���
�')\5fŋQk���M�r���b�'�~-2�+��'4���Ůe9����'��1gOJ)'}.��a��^�F�'W�1�( a��IJ�s�ź�'"D8"�J�,�^P�"�ب@	�'�ʀ�F�9Q�  �����X��'�p�Z�-3�����5{?���'���-c9@yq�U�i���s�'�5��A�g*f�)A��$u���*�'В}�%�G(}b`�e!Эe���Q�'�Xi���2���@�T�^x�a
�'�^dk�D��h�J�Q��B�d�H��	�'o���� ̗Q�l��@R�]� ���'ƶ�3�ʑ�����F`[�J���'��� !L�,Dl�F��6}� ���'�8#R�F!*(@��5CA	z�����'Ϙ�q� ]�h�P�g�fMT���� �ኃ)4�J&ךF�0�x�"O�\��]-|�9���G��0��"OTE�2cQ~B(�b��)��"OD)@p�1�uKЧ{�a� "O؈+1��6$\�s
�<4�d5h��'��I����I���˟��	���ɮv��U�d�H2�4yQV���Y������P�Iџ|�I��<���� �	ğ��	1A�p��	����kL�2�
�������IΟ��������Ο���ٟ��I;1�.��K
+b�`� ����QVD��ʟ��	̟l�	��������	ş4�I�E��z1c&
ed�01�Ř{�D��I��Iџ����� ���� �Iڟ��ɰ_��չ`H���z���Q*����ڟ��Ꞔ������	���˟��	KwD RdL�5xv�@�2��KJ���ퟬ���d�	����	�����ş��I�2��`���!/'�Y�!�GA:\�Iʟh��ןH�	ğ��I�L�Iǟt��	G�<�c�Z33�I
4ꉲ�d��ǟ��Iڟ<����h��Ο��	�L�IN�R��B�a�0��A����-�I�����	�p�	ßH�	ӟ��%��h	�+[*������ơ:8|�IٟP�	ן�	������D�I�$�ɚ'���R�P�EB�D�w��*���	��p����I��t��՟�I� ��5<� ��QgҞ�ꥂF�՝a�����ԟ�������ϟ\�I�X�޴�?��H����%#{�$h+𨅮ZH
��Z�H��cy���OڝyC��<�&prQ�I;�D�xJ�|V�=�3�� �ٴ�?�v��j��<�����8W���Ye�Z�cV(��ܰ�y�xɢ`�9"<l�˭����,3c�t+dӘ�͓paT9ч��4|2���ӈ��	�,e�I�<��oL$?#���(O��' U��']�P�P��F�R-�C��M�^��gLțe*n��<���T�F(�'��7=視#C�!J��<tH��j����O��Dγw%�1���/'��?yk��PѺ#U� /s�q�*��D�D�O��Y��'���jTΟ�yS��dd�,����a����1Y( �pef�<l]��[3
�2���INyr�|RGP�<Ȉ9�yB�ڦh�����E�>�b��	�m��k����dZ}��'�)ƚ>����WBz�E��H�!!Z��+�.�@Mȵ��B��yb�x�~�YA�9�`]>��QG�OZTÓ.U
`$�HqR�L=c8H�R���
.O��DN\�v����9Otʓ&�D�)�7L�4���j�(mu�@͓����g~��c�d��Ц�1��(�v�ە_���A���lL���Iτ���A�O0y�	�.Pzם= jh�
��fR��S6m�!KrlQ��ȅ ��!�'��pNn
Ư�<�'.�rw�ݐwU��Q�d��!��`���0<ꚰ)��Pe�R�'4���K�՘'y��A����թ/TF)2@�>]`h;�ǸO��' �'-��+è�O�UB�/�-��)�� ��R�Ϝ};ƴj�C�g�x�R�ޯ-�.���i�|؂b�/^�������?�$�#{|�
�
��-��b#�56~�"��,l�˓���'�$��|yW9OLP��D|�QT�ϻx�@�6O`�m��H �n"?��<���?�A�S-�G�0X�pM*��Z�2/$u-y�>\��i�:zr�����M3�i�M�i�	��Dj݉2���u���7,��a҆��	]�,�z��P��@q���<��S��l?�s���`"��rb@�q�x��ٵ�,�In-����??�b�iT�\�y��������=_bBy և��x����O��g
,;=�O$ʩ�V��6 ��j~�X�ٴ<�4��GC"bХ{S���P����o�O2Ĉ�i�Ny�0O��"C�����?�5A�Ba��b�ۦ}��yjcɓ�<)L>	����tB���<a��Pl�G6P
Niۦ�C$�����&@a~�O�>����?���ɿ|P�F�8�8"��C+��ڧ-� �N��Wá/C8�A��iAld�a/�)I96<�'��Έ�XrJK��˓\^��bSk�.��g�X�6,���'��ĉ#�y����T�'�\�H��d��!1HĢ��4U�f�3�;��X�3�G�@��*�M���=3���'���:�&�ʁJY�a{퓩IN�����F��6��[�蹹�(wAP UF=��D
f��eR]w>��0���<��.R�V�(�d���Ș�g��џ�� ����l0�?q���?��' ͖Q:.���v��j���2!H\�1��Dp�iH�R�bh
_*2�'l��O��q��m���M�;c����#�M+�Ǳ;�� 2ði��6���䂄H��̟���qݕ�ק??"���͇?�k��L%�a��,���C�O2��$�`y��O�bC*��)��dT"JԔ�ES+-�|��+U�;�"�$�OP���O2˓
I(�r�f ���$�OT8��!͐�R�#��q���O���D�On�m��M3�(�Z?���Q�.E@�r�R:��ѐҢ{�*`G+�ҟ���ً``ɹ���<�Iغ�����u���J��)�A�{�=��O�j�i�'��'gv�IU�Q�@��OU��'��۰\^�}�S��*Z4�ؔ�V�I2A��K�,A0��'2�z�$�D��8��i�`ӵi��+���!ŢUAD1nq��@!E��M�2ƢI��4�Yw>�ȩ3j�O�X�Ȑ��u7ʆ	�t1�Ϧn�T�p&���<橛P��ky�-�O�%�@AB����$�O��d�V�je'Ԛs�n�(vA�>)_��Aq�(�.�G�cT���?����?)�'_t�Aϧ�?i�&�0R��ۆ�qE6ۡ�Ǯg�ɦ�MŴi:TI�'̞�AU����)W$q���V��E���53�!�F�k=� ȋb󄍼M��I�����|
7_�( ��XR {�N1�n��LM*�,X�w��&W2�ϓ�?9���?y����d�9zU����O� �t�ýز�ChW��t��V��Of�oz�Mk�@�V~�>i�i�̶Bf� l�Xu� �wݶ��s	��%n�Kc�*L*}qR�
0?��Y�!�=4�PE��JF&(�E��|����� j��m�3���W�z?uɂd#>�,C��O�$�O�IƁ)��.L�c���s��J:7�N�P�`R���O��$;=-��#�<��i����&�~2���'�Z�7�ɶ\��N� �xe�5�(��
D-�Mϧ{(�urXwE�qJ�<O�H�oR�1|4�
�	��8s� H3�
�{��*H�S��h���5����?���?�j�o���jӏ�U���3��ɤ�?9����D�97����O����O@��&%��K�6tT�3�"?#��YZ�� j/O*��vӠ�z��OB�I�ą����ǂ3c�X��SCql3��^Z{�Y;a��p4��Eצ�y���	�Px*O�����1@mbT�ƚrh��ˣF�֟�(fO(U ������ßl�	Ty�"�hD(p�JH�|�I��P��Ip��'_V���O�0n��h�D�#?!BX�ln��d��)t�<P̈́�Z��b�ƕS޴#�P\ ��W�#�f�4�$�?���w���'{��B�7Or�Ktd��p�t}�����j����U�>n$z�k��?q��?i�'zj�(��`�WNU7s�@rq��74��pf-DB��	��<�����bjA�|��웞w�V|�	��.m"���TS��K�e��LoZI!��I_\A�?E��F�w�����ɇ�W�JX�"@P>}Z}P�e܌�I�����'6-1%�<t�'�����ҢF�C�m �`@��%eJM�t�ĥW��'���'�	�*��}:.�Vy�'�0}0w�>ո$�A0Pny��Ȗ����B*?�W��ڴ*���l��~����LC ���(�(m�"��}�l�d�G�<�2���1�!ӗoC�EZ���O��p��������M���;��ʁml��J0ȷh?����O����Q��,;#�(�I�O����O\P[wG u��Ѐ����s�I�O���  U�i�d�Opo�џ��s)?�;3��UVGZ�4��<�eTs
2��A�(
�z�i��y(�EVHd��f$Ai��R��$��Bܘ�jEi�AP4e��aނf�F5q2 L9�l���	Z��-��'�B�'u�4�UQn���al�{�`�t*�`���XrU�4� a�2o4�ɗ'���O�6(i�OVR-�#f���7@M/��٪K6F�r�1n���x�r� ��O>a�Tk�.	���O��8���g��
�0y`bT`v��>/2�Ѥ��3�yrFU����5k�3/O�%�	�jP�3)���9�=<fN���C�g� ��џ0�	�P��wy�
?L��}Pu�'
�$����$ ���eN��i��,���'�H7-�O��)Ř�Tc-O���j�@����N&���sj�1r�Г����N\H�eɧ"�X�����O��+����u��
���ϓ�u7���IJB�H�	e�	B�O�� *��A��*`�OP���Ol����<�b���T�F�Фe5m��$��"Z�TN��O���G�^�xi��<	ǽi?RⓈ�ybJ6J���C��A��G����,��'_�(��͊2�OB�Mh�c�%K�Q��'��a�G0F�ꨠ��Q�DOhY���P v4�Ɍ���+O� �I�V��e�"cHݟ���̟��鞿29h�cM�doT-q@+����^yr@��cf�1t�'|�'J�ԧ�#�J�Id����Ik2$Z�*�h�O��'�"6mWȦ�xЈ��@��M ^�I��;��8�B�3?���h�
�,�ʡ{#���N��4;ä�9rP��Ol0��?7Xd8�_�L��Ő�R08ss��b�v���a��?��d��*�tI0���?�'�?q����GV��0��e�Z^X)��MӚ^i4���QS�����Oh�m�ǟ�3r�6?��V�mZ�`|z��V{(V���,m6ЀݴK�E�g�̉!�|(��a��<�D��7�H��V�*50O����\�`V���ࡁ�MJ*�A�'���X5OdH�-�O��$�O��	ƢEZ�'h@4M�c�׮@��DX!�ہtaƼ��f��n���?)����D�C�|B��ei��w7|���O�x+�#�J w��A�q�wӸ�l�A$��ɣGs� ��?�5c� o8���&f�XDQ-� j)�t{�A�de�牕F�U�V�'���A&��<���'��WgǏ,�r�-e�$�J��ʷ2�2�r��ϋ__"�'b��' �3�<:��A~y2�'D������3�l`�*ʘVe��%�'�f��O��'0`7�Kͦ��O�����o�? �d��䈐?�v�PW*�.4��H�5Omq�����M�g�#E��˧��	'�Ę��
�D�V}�T!�f��H`�Z�n��'"��2~�M�D��D�'6��'��-BSm@<-�(�SDe�Ա��'�^�X��~FB�'��7-�O��D��杻H�R�`��ؽvO��s�e��/氹kfBI���\qߴM���G\6r�1b�Q�<�G��+[��]$M��!x�IU�4	�80��M�88��N�dyb�O�u�w#ж	$�$�O���r!`nU	OF�04O*jNP�fk%<.��tz��;�?����?���Uw$��'�?ɷ.Šb 4+E�	��#�0�6^����4t��f���~��mj0X����:�K4,��aa�\�/�����U�L��t��o��x٢��n�{ԉ�O���E��ky��O����NV9(Bz�B��'��/�FM��(�1�y��'�b�'�X��qf p_ ���h�h1�׃2^�A�g.ҩ1���	��MK�,L�q�'*Z�\O�vl�t�Pt�'7Ȍ��mּB�Va�e��d�1P ͽ��L��K�O��� �&�ug�)\��!��u7���<LX4"��~��y����U��X�F�]&_$��m�O�$�ON�II�!ʀ���.V3�2��ʙ�]�8h
DL��d��O��D��~�,Lr�%�<a�iP�c �yүA�`6��b/E�1+,���J���'&ҼH���!T���OF`��Ec�$���'��t ��!�J����B9LJ*�K6�xh��>��U�.O���I�f�$(Sv�Cܟ(��ҟ��/>��Ƞǂ_\�j��PKG��L��Cy�Æ~u�9��'
R�'z��͛�g�>l���t0p �E�K��3�O�@�'���i:|��'��ؓ�!��|�k��*�� ��X�V����XF�`pɔr�eL�<�2�T��2ln�'7�2�@�#�\��R۸Y�� �O(��ꎱR�����O��O���<��
�:׼4�R�f{�:�8@��/�bU���Z#�?���̛�'��L��O�'��6ۺ.Ӣ�[�a�4l (���2?F��o:uP�<�,@�{Ĵ�(�/��x��J95d��^7-��{��� z����O4.D�"�q5���'���dХg���Z��O�D�O6���*J_��'4�ʵb��=\)�l���9&�."�)Ǿ
h�����?���ڵ.V�|��7���wv ���B([�h4�ׄZ�j	TA�dapӘ�m�p�	�"�Э��?�#woT�U�lT���!|�ܛs�J�rX�18�cW����	<4�P9	G�' ���6��<���'!:�AR��l��f��-��&ߞp��9iC%�-4��'6��'	�	�p �A� ��0�	Ο�3gJ g0��;Q�6�����	���Cg%?	�]���	ʦ�y�nF8�?�Uς*G�&E3��ω= ơ1e�>{W%��#4D��Ё�r،;��ֱE��O�=�fݽ+,BQ�p�<!��Ѫ1GφK������t|p���O���&\h�UIU�'�	�O����O��"��v���W�wW(ѷn�OF0s�n[��v�a}��' �	�O�.��P��U�K�,���������urĂ-@�2=nڦX������۾5�B8����)GTn+�E�4>�����a�>� U�0">)�p�T')"8D���TM}���OrM���3X�����O�D��.��F�"��e_7\��1!)��(�ʓ[�=�a�@��?����?��'FB�	(O��3'� ���Q�Q�Q�*|N��£O}��pӞ�l�V��	�,�H�D�?e��@ň����2x�PΎ�eX쨄.�W?Q�wMk����Ŋ@��e9f�>q@'�OD �w�S4/,��%썳��v����f[�[���$�O
���O:��<I�E(�����w*�Y�Aշ�* ���d�e͓2�V�'h�x�O�t�'��7-	���S����~J���cuRy�V�K3U��3q�JcZl�z֮s�,CggH���R�@��'�V�5�w!�`�w([>Bne�4�A�5W\l�PJōG��Q��'|"�'n�4�Y
!��y׬��
��E��<?���M�*
���'\b���}MVu��\�ȑݴ�?����<a��97pX�f	�/
^L
���'T�t���LVF�K���M��'>��hv	̨-�z�	�U_����.�1"'�Y�S���5�f͹��K�*��I��Γi:�ȫ���ʉ��.Y��?����?1*�}M���O5=Ε���?����K)�$CÍ�O,���O$���){&D��D�bBb���N�-(k%��L�O�1oڴ�M�f?�u����������(���70Z�a0b����Y�/3V'�$3Ę'I���	-��{��'Z�}#��y�@��+����ЇL�{y�	��B4H;*p��%7|e�a��|�i>��I���'��9��G(c�nK7c�VU��H 	��V��4�?9c��C~n�<y۴i�$C�L�>�ReЗ
�A��رd�i�u�C��@�S������d��>_P����,=	0	g� �`�ف$B��A��0���Y��p�C�OJ�9Q�C1L0V�D�O���������̤|
%]8k?��a�qM��ŋ��vf( `q���On�D��ę�EG�<�D��y���%4���%[�5@���աW4)���$oӾd;��O�Ls�ب$��O�b`IT�W�{_�<�t�d�����%�!;&�,�g�P��y2K�x�,��4W����'�FP���'_ȝb��IdҀӣa�qQ��Q< ��i��$@"�'fb�';�|���I�d���	ӟd�cC=���aM�o�^5J�Bǟ�*!n/?yX���4<2�f�ۉ�~�bןX��P�dǃ�w�T�b�T1Qє9�4�]�<I程�c����mz�Em��<Y�M�p���D�:GK���%�KL|��`�B�H%Sag����4�?���`exrd9��'�?Q��?A�.@-`	�Qa&.F~�`�	BY0�?QT�:u�hy�/O�o��AQk#?�;r�����0J���ᘅu_ܠ"ǨH���Qt�i|6 ��ڀZ��-"��W��y���,ȸ��;v�h  ���9k�^͛צ�v��$�RR�&��5ym�%���,� 鷌��l�	ӟ��S"8��v��l���n�N��G�H���D_�h�`5¢ �Od�D�Ob��`i��,�!��%��CJ]`���	#�|�@R���46=�&�3�~�k��[i։�������
/ �h�pࠒ3�:�i���8㪔u�D��yOքy����	�r�	�'�fM`��'䞕c�o�e���ƨ�*�$��g)O�3�Z C��'�2�'���'��7(J���oZ��8kT/_  U�q���ԋS�rQ�j��@ش�?"�GQ~� �<����MKֈJ�T��k`�'S�l:C���v�BI�CZ�,�X�l
�=�vY�"�[��[У�v������\�RYi��hi`1�㛩@�n�c�.�֜��.�;'�M����?��R���{'-�,B0$��gl"w����թ�?9��?9�W�jsĭy/O�9o��\��f���Eħt�ԉK�(�	�n	��K�98�����?�� ����Ǧ��7<nV�C��ڣR	��9)=F4�`j��܌J�N��j�(�3�gݕ	�b�:3	,�I�y(L���NQ��C���ş���ӟ�qQ�ݞ��| ������ C�ӟ���Oy��� Bb�DRF�':��'�����-%� �
W��`��HK^��/� ���z}�Gh�~Ln�(wZ���5Uu�4�����L�����L���ҡK�h�ڍ�.��	��!&iI�u�A�3O��sO��?��R,s�����<Q��g������Ǝ��J�2���O&l�3�l���O���O��Ģ<��cߌL�����	!�i�!��5$��Iv����D�ʦ1�I#c�H�"�	��)��^�l�� QPLuSq�֑�MC�kM�Ε�@�������2�(2+w�U�q�ܭ5���1MZ��$�!v�b�K�2/t�T.�O�=÷K�R��$�Oh�D��N��a(�|��>p��U ȴ����&[
�>}SG Ū�?Q���?��'c6p�	-O��mz޽�p�B�d����V�.]���s���MKռi��\*�'HRH��6�z��Y����]<�X!  ���Q߫+�^�Pk�<���M����DՒ ~�S6n|��I�i����H͟0�'n�~�d��g/O�C�θ��K��� �Iǟ��IByB�"#;����'b�'B�{�� �zѲ��]�2��4�?�Db\@~�g�>��imp7���=o���)u��d�P,}��	`�"�6+MX�� ��H�cଲ¦ŌT3ލۘ'Ք	��'N���'��,$�D�L�<��z��w�f1z�'���'����Lכ��O'r�'�BM�-|��8PFc���q�NP�����@�D_����4�?Q`��B~�wkH	��oM�]��Y&�
�E�Nl0��[*M�xyCfy��TICN��Ւ�PM�)�DN��ԙ�Xw��� ����ӋRRM� %My��Q���s���:�$L3�h!	�,�O@�D�O��iտP9 �f+�f�*T�L�.W�S�L�<ɒ��(#��b���?A��J0��0��D̨9�����T9j% �H�d�D����'&�7�Ȧр1鵟|!���<J���`C�CS�-����ʙ~��h���u�rQ��d��D�`��Tk��-H��q2O�5
��O k������+�¢+^�R`�K-`�t��I�Op��O����O��~���%�ߊ�y�n.rt�d)�.m�N �`��<�g�i��(O�����Ky��'�&L˸.QrIk��W	$lzհ��	?�0@Э�rʠ�P�Up��OpQ�;2���R�j�����ߩS�G�l���!1c�T ��w�RT'P�ɕ��ן(�	�S�?�TP%?�]M{fu2�9KZ&Y��C�:����柠�I�~:�9�u	_^yb�s�4��n3&牿Ye���D�(;=рY�LF`�Ձ��`��Ǵj^>tnZ�?��7\6(;L|��[Ο�C A���l@�˘�& ����ډpQ�'��z`"�<�@�'yrpA"��y�2�'8�byh1�"�Ԭ9r,ݩ /̏CR�'}副&��ۇ�l����ޟ���6W8�!n�-XpU2���#ez���!?��\�`��̦�kȭ�?	 H'�*�X�l�f���&�<�bA�L���T&< c¯T����韒�`��'�vDđ�ذ��݉4",���(�$��<A�NX��?q�N �w[ҨH��?�'�?�����DS�7�L��'މ�~�h��B2��̀��۠��ɏ�M���:�^Q�'j�*��ǝO�2h`�&�o/^�1��^�R�7M�McL*2�.+� `��O�}:#f	�u���*�A>O<$ғg�\⨉�)9P�����'����V�n����M�OJ�$�O��	�z��'A��z�dP
V��1�A�z�h�qb̟:�\���?����Bwi�P~by���o�ּ��+�I��I�'`�mڂ�McC��>aB��-�zq�ON��$�Q��ؓ嬛T�҅�eN��h0��A��y��� �\���+B!AA/O|��	�)���B�N���r�f�e�$����2=T�(��	័����@�	\y�Ɯ�a]����O�$�
(�<���̉�K�8K��$K�0��	-��$O�����46ĺУ��'�"4�/%j� UV� 'v�4���!?J�8,s�M�uc�	�\�$��<�\wc�x��0Y$A�2��$*�9��M�9�����n�"\6����OF�D�l>�!pǄ �i�O��OR\b�m�<m�.UX�Ա`�"U1u�Oy���Y�LFD˓��v�'>����O�Μr���4nB����!�	bb�!��f �t�&=lZ89Pl�k@ �/�j��g!g��K�㖳.���K�~�F1�`�YH6,;C�^&X���ш_,��ԟ����������ݟ4���?E�+�']Z�;[I"�*�l	?< 5�AZ��1���<�R�	蟸���?��i(?�.C/r��U��K [j�@MO��WҦ�[۴ �� ΓG]����스���'�*�� �Dm\�14��M��HL��F@q�
U�<yçS�����RS���'�\���*rd��
ٿrh���@�����S��@V���O���Or�$�<iN�7a�Q����	�'øY��t���:��<���?����Q��|�,O�<l�M����d�YХX'���
� P34H3H�*�0��Í��?�D��4�h��c��	sA\\ϓ�u�B��bP�4�ai��%;/8��שK�)��@�@��"�'�b�OQv������'�Q�TkM�*� x�E�V�O`�lR�'���'P0=)�����$�O��䐅6��ȏT0HcC&�{�@�
"ш�X�3O�� ����SŤem�?Ѱ�D �2�&���j�� �T,�g��F�l�Z���ݷRվy �'l��B��<��'�F��'n��(��'�/�"�VA ����b��CC����'��	̨܂���y��'<�d@��F�4���@��@@],a��Ox8�'7mX�AqA���$*,�7j���� ��g�P�?�r����A�JèmiAǑRRQӳ�,J�dzݽad�O��ඌ�@y�W�2��Щ֔(b`xC�ʅ1:���3H�U�Q(�O��4�����Oʓx%<���.ӕk�z�Kt� �<A�ԣ��[J��'
7��O��yВ��h�O�mZ'f9�r��U�}�0}гHN�� \y޴{�L3r��643Јʭ�?y����Y�(ם��"��u>O6��f���pa�fJ#Q�A��'V���R%��>pS��'|��O�e�1Q>� o�[H:����$h0,	����N<s��t�L��П0�Ӄ�R�4���wU��Q�0��(bc
u��$�Tiq�J]n�2�Đ�P�V�5a�?��S#{�!�H�|��#R6/e��6l���Vy�@�!��6n4�$��M��ʓD�.
'X#tmA��'\uH�gN�V���rA'<w��%;t�'U��'_bY�d��jڸ�t���8�I�6����mݬE,��r�%j4�I����'B�I��M���ih��)�'K.�,�fr��!��5M��E{�����|̓kRY��˘5x�Ps���\���/�?���"R
�U+��7����&�і\��( ��O$���O:��ʌа��v���O���ˑ3s��CՂ� r���P�x���ֲs�������O���Ӧ���=s� �Ӽ������:���*�����c���!���c�\��xY?�X��f�ɟ(H�(�1k��F�-F��X����.b��1��*D:�T���V�X�I[a�L��?	���?!���K�Hā����Aݼ9���`
$����b�ҝ��,�O����O��IM/x��ӭӆ�!�d|��nRy!$Tz�O�!o��M32O \?�ꟷz����S�?id�يX$։(Mç�t�ZSL��"`�E�Q�6R��,y�p �1O� ��<Q��'0���!)��M"�D�^��e1�C�'08jB�'vB�'�'��	&u�2tˡ�Pşx8��Ʈ4V�q�>�B� c�@
۴�?�G��`~"+�>�T�iJJ6��;��9��k�����T���}HIˇ��&�>a��˝~���D��=�[w��ȓ���<9_w����s[B ���!]�R��R���j��
�%$Z��D�O��� �2�9�9���[xr$0:�R�X�J�j �O��d�O���́�Pƈ�����'"����'j�ZgM��W��ȥ`��I�^��Ǝ�~"mٟen� 9����b "I����iH��y�&���� $T� #�SB��dJ_=bu������y������I��?��Ѩ,�s��?����౥�X�R�<zW�˿3�8����?�,OVP����:�@��?�'���+�L1����h��-�Pqcj�z~�Ͱ>qu�i%�6-̅fo��ԁM̾�Q�O�T��udӁ:"� W�O��i�/\�x�����O؄q�'���Ȱ��#�$	\˓\��`!n#(�@p1e��?f ����'�毄,j����D�'�_�Ps5
�)q�vLRV��� ��) �=t@�C�]dy��a����R#*��ɚ������:�E�CJ��{Q��_���R,ٞ�M�PԦb$�-�b%P�7�2��,�i�bz�]!�Q"��ֱr�Դ�%�J�*�4r�-WV�b��O� �i�)�^�D�O��$�8s�ʲ|Z��$f�`��3�W�ڵs◱C`0S��?����?a�'V�r��+OX�lz�9A�hۉy��6A��=��50eD���M;"�i%����'�������2�'P8Ūq�ȅ.f��T@R=���� E�\��A�"#��<��lŴSx�$�
U���',�dȜmn(�zF"�Oj�e��J�y�V��~S6� ���Of���O4�d�<����o�2�,O�d�+I��J� ާyP�PQ�F/R�D����������ۦE��4"V���aG�y�"���X�!m� j��I�b(Y�%�~�	K�t���*��Eaq�d�l�;b ���!6���GΜ)��CF&�-=�l
KI.W��'\��,a��hkb����'��wܔ����$a�Ԙ�,�Y)T�aW�',P�	D�-��ğ��	�R_��Ӽ�1O�8Q�󌌔C"��a_3PY�'L�Ưf�;������0C����'��S�����#;jhX��+7*�xm��㑑:-��kE!�<��'�L�/`f���'���'���ڕo��u���.`PLQ��<:�h�H�]�� `��Q�����X�	�?�Q�B-?a �� �����¿W����4`���	��M{��i��Q�"�O�Yjv�T���V�V�x��cM��B��t��Oۚlܩis� �,� p�?O���&ɕ��?�3'��u��I�?Q�+�8S|�b�cG�T���nWZ�&�0�)\��?���?���?�+O0�d��i��DI�2(�l�E!	�\��M��E2&+�D�Ԧ5��6X���([����M��iAN��`ީ$H���p֟V��2"�����@'6z%�M'�'Ofu������ώ����Ѻ�@~��4A�(q��/Ʌv�X���.��2�z�
7�����������|�&?�ݶGM�8H�넳g�J=r��
���	�	�6��**?aw�iC�Y.�y«�b�*��r�ͪa(�yC����U�+H�(��
*!�+"�h���I/(T�Ye&^�q����>�6@�G6�(3B�Qq[Fi�?	`����ɚ�?ap�]C%�`���?Y�k�>��tGU�B�6�0��o̥��?�.O��e���(��$�O��d��ደl@�,�xH� �G����ኻp�����D�O�7�$�<���h�U[BJ�(���=��׊.cT�����,QR��s��-y�>�	r	�<�Zw�r��d3�W��X�d�:,'P�%��S�hX�
D��?���Xu�`��O��4�p���OPʓ3fx�B�ǲc�N��$K�E�V@P�*[�4�����?չic���DPe}�r��e����r� ��l@� L�4���]+B��M��pU�զ=>P�	8�d,I@��^�rC�߶�y�gZ:m!`���A�;t t����?)!�'���	 V��'��O'hp�gQ>]"�aG�d��-���Z�Z��a���64�8yc�&���I��L�S�;����������U`ܱ���6���h]����(� �Vi{Ӷ�y��Op�p��e�d�O1��e�QemT��� �rі�Y��)mgԨ�G��yB-Q/᲌�ֶi�f�:�T�,�'5b\���?I��$	RDs��ԬE ,$���?����?�����K	O<��4O��D�OB<( ��+z�8��7���̀C��O\1�%��P�'n6��ܦ�P�a�|��IϤg�Ȁ�ɇLh��#&��gm��4��؟ Т��>a��s^и��'~�4���yΓUgr��� ����:�"i��Q��M������Il��@a��H�؟`�i��Ç�(w�Pf$
,
�X�3oӟ�6���Ȗ'g�6��O�\ᜟ��'7���c�'Zw~-[��94p
]�*��~�6��4Bɺ-�RdƧ
On��2�[+�?yf*�}i�֝��AP+[v�iۄ"��f-Ұ��>f�ɵ�?a��G!|�Pj���?���Z N[�\�l"�Մe��1r�e�}+���?��$2z��ڧ��?��b\̉3OJN~�@W�j%`4��!��2��M`��ܕ �r�'�T6mN��)�k<"�T����RЦy���u�� &3H�#��7	�)p��ԮK�����%�@��'c��@H"BJ�V�����D@ß��B����;�O��#X����l^$�T���b�,��ޟ��I�"ҘE�'70m��+Vf���GT�[kJ(�5��#]4$�[���Q}�'��E7�y�Ob�I��M�ѳiw@e�0A�J~�0��A�e������|��-p�5"�6�#��'zΤ�W����+��"�y2��TXc$�P�� ~�$%��D�V��(�����$�V���'y��'�d�Xo���y�EXRL��+\�_�(�I�q�z���'�RK� d��s�'\��'���\5�y"n
��fY���3Z�e��J�z�RHv����擙w{,Lm��?e��MY1v�"d�х�֟����3�b��O�2����T�" ��'*����<���'�U��'k#��'��'E������aB�Tc5�@�>A�1�Ƀ�V��'���?���ҟ,�S`������,]�����g	�&���q���I^y�EoӢ�oZ.\.�۴[	�ղ��;���kFQ�zQŞ�/�*� P�aӜ!��Mв4T�]�'c��<Y^w��ts�{��U�W�$i�M�,cR�X�J�nȒp�#!Қ�?I1�O4+	� ���?�E��?�fO���$�<T܉!�����x���W ��%�[&�V1x�j첆��O�XiA�?��ݴ�?�W�i��A�A�4�X{+?��p��(8�������则�'.b��3}���R�l��M��Q�:O�4%$�!H5ndy��ŸztN!�W�'����@)Z� ��O��$�O�i��! ��O�u��*�;��b������@�;P�8��U�i�*�$�O �J#ʨ���d�8�I�>C�YQt��<{�d@@�)HrE��4[��槞�����1�#>٥�OY�ם�;���$�E�C��� ��%h�7}�ܰzs�'F�z=��'���9���?y%�קm��w(�F�6����S�'�ƨ�U��"?�� ���cB�)B��'Z�'	D���W�X S�@�y/Z���ޟX�	���St)K�w��Da�[������T�П4�'�6����%��MQ�M�嚢K��2H�Y�T Tb�$�4��?��#υH�7�ˮ��u�.� l ������e���-L���/sb�:Ɔ��?����?ɐ�:O��U���?A�Hʿ�?�ǃ��?�pI����x��M�Idl�bfC4�?��	#���'�д�C�'4��'p"�'(M2$͜&p(�Р@��~gs�j��p0`��b�f`ᖬ�"��T�4�O�9��A��B<B�%X��)PG�'vJ4��Q>R�X��̏�\��	8�?���?Ő�����?����_������Q�?Ĥ�RG��>x�y(/Of�XU�A
	,�ʓ�?���_{,�O��L���G��S]�����@���Ɉ�M;�i�:e{�'�4ikW`��J�'w�H�'D�of�(1��)=����jֿ\C�`i� ��<�)�~�D�;&��m�'����.[���#Fݽ1HV|:��Z"���P)����O$�d�O���<�V���������iR�Q�0����Yzyϓ7��F�'�*�O�T�'Ѡ6MEצ� ̧&>b%�ҩ�-.E��"�K$C�`	G_�3������Z����E�/'2�Ό*?%�|��'`����u[���u �)�C33
j	��,���Y��KΟ\�	џ�ӈd�x�$?��ht�a���
v����eˡ|�j��	ߟ���b;`CMy��|Ӛ�DJ�m�Y
Q?4D� ǅ0B�<����K���(��O�m��*
�6m�j�ʷf�0�r����O�ͫ棛�p����G�@�sP�-�Uƅws��k�u��4 P�0��#~�1R�X��?����?�1�_�=]8����N��C��7�?�������j���Q6��<���*�`��XOj���	W%���K.�Bԉ�'h��?Y�4=����}� ��?qӔŜ�7��rJ�4:����&g %C.��rǤò*��\�kx�H�����ɩGV4�9/O̅R��@�yI��1��F=c�D؄(��f^'h��Iҟ�������my������&��*D�yh4"]�
`q媏-'��I��M3�b����'/���M� ��$�@Q�� S r��R��F��$�W��ȗ.�P(�X��'Jt$x�@���Ó"A�_ݎ�I/T��bѵG*��Η'bp��^��21�̭].��	�L���?�j��H���X�5^����$Az�DٖÈ��I��L<pK��'02�O% �*�O|��i��n7B,��k2��2�Z�����Xнi{�7�B��D )<���˟&iZ�
�3�|��	W�( vB̰:���S�M��D�-����'��xR�����9���Ғ���?��_�FI��׹�T�+�m��?����?A���ڋb�yiׄ�O��D�O�l��6}���7��6�`Y�d�O̔�U��H�OL�l�+�Mk ��T?����e�N�l8)�E{��,8�^���k��;�c��nv����J']&�'�4��E�8��C9)2���+!�� D|2�'��LʺP�i������'��'���V
!&���sɊ
 5���'���c��,p��'��7-�O�����]$(�0��3J0v,p���2��D��/�_�ڀk�4��R����aQb��#��<i0�ՠi��}�I"%�30OP�C�V=mX��@I٪vN�^�(���B��x`�!	�?����?A�'|�r�2K�RE�L�~l��LN&���;K�T9Vį<!���£
@�|���<�H����9�T}q��9Qv���b]���I����㩽�X+�ǉ.������CIƬ%�$H���S=LELM���D_��Z� pM�ΓQLȍX���M���Y��[㟜���J�n���GMA�G�| ���,�X���ҟ��	&�}�	�o@0ݕ'�>�)����$��#�,��lO;.����!]r��U#�5�"ρ�y�O��6��Od4l��MKELZ�\��#�kE�3",���F�^̥�G�֥Up�)Cg��?a�`����gˍ �V�̓�ugM���Q��,�����k�"�*��mȤʂ�X7�?���?A��=�ji9N~λ�.ZW#1j�4]�QFؙ��@Z��?��>I|�M	�|B�{����'ȭ�'���c�Ϥo*DmB�'ï���ca	��~R)ү*q�Xռ��4�ؾKFmj�(I(�yb�N;?��вʏ�A���UnZ� +<P ��<a�ʈ������2�a�7Y�*���؟h�I�_���M�Bx�BB�� 5�d!�	��'O�+��y�'�B�O2�hqul��!D( ��▥ p���)����o}�ip��m�EB5��G��m���e>��fQ)62�X��)�>i<��.^�=H
�[��x�D|����#����o7�˓E�%��'�&������q�����'Y�,Oȿl�����$�'�"Y�dF�+�U��ʞ־���/�1-O�-�$��Ey��bӞ��C�5��/���Ϧ�J�Ԯ'��4sGh%j���T�M�M�Մ�e ��2 L-T�(Tϓ\F�q�q�	��� �S���K���Q	�37�`�SnݶZ����O��Y��M������O��d����x!�|��'�%Qe6i�v�M�#�Z���$Th<�I\��?��?��''�j��.O|�nz�b�ϖ2h��;Q�46ռQ�Ɔψ�M�g�i�J���'�rI�q���
��h��b��M6{����F`�
Vep�1���w�F9�I��<Q��	 ���D>Ғ��'J�$�W��l#��OfT�פ�/���	����a?�q�'�O���O��$�<q�A.&Sz8���?��w��R�d>��|)DK#	-�l0���z�'0J�E՛��y����OV��2�\�b�E����	�u�A�3 b�p�( �I�Kf�p�"_�oC�ʧYa(��ɌSTx��tƔ�?��qJ@�M�|��!P�0SR�'��'�O,`y(֓��'b�'���;re��d�����FnN�:$�'ްB#M͘/��'��6m�O�h�4����6.�|j��!v�|2�#�`��m�A�� *U�k�4N��	r��@]`�Df��<�$���v�}�}����A,2吖�,)���H�J�-P��'O��$��T��p�Ri�O���O4�I�k�R�)V!Z�.ʘ��`+/%��Ɓ�<�D��a�y��?������+���=Dj�5�Q��#2����_����'�7�����q�����TD�:u�%l�8� �db��S0(�Ă�l��4� [C� �d�ؽ�>O((��J��?a��Ts��Ʉ�?Y��L ��dSQ-6^��)+�'�?Am�H��^��?y���?���?a+O�Q��J��{L��X&.�����,�Q��A�珇�%7����I�[y��%��	��mڰM�t� r��J�(I�H�#~�CC.F3lf�XTAQ�0�T���'�`�(��A8à��y�������4� �&�H+:�,���!d�:ؓ�'Y:8�������?-#Y~�s�I�:�v1ƥ	�FBP���Kԟ���ӟ��ς5r׶H�'e�7�O�xAB0Oh����)8�:"��/������ L��D�&'\�j��p���ɋY���M����R05@��=0@#7�7|TR�͆.(����D�W��'E��$E"i�\qJ�`�O��d�O�Ts��\
��y��Ƶ<��`c���O��d�<iA��z���Γ�?����j�G�Ne�D��*v��I@Ff/y0���'���94��!l�V,K�������K�^���6"Թr��$r��ڒ� �6$�4��}��L:
���Db�u����O��Q�'"�� �@X8Q�D���O�7��1x�,�O�%����0(��$�O���OD���<�����s��Ȼ�"Q�ީ�"�Q�v����p}�	�M+�`*���'^�p.�f`�.@�{�C�#$���� `Â)9�6M�(i@j� t�X
{�Q���OX�y�/�u��ڄ����|nd��@�E%x�-!���5p�����?���ɪb�(���?a���������G,C�TuQ!�ș$5b$���+P/�t���� ���O����$�"ԙ��;�����[�|�����Ĕ�-�2��Q����}�(4�k��p��F|}����*��f�;,�rY�7'?2*$��e��H����	<�d��N��9��Y$p��R�x��%�\]�a��?!�LM-��i �F�XP���?���?�����J�p��ۓ �O����Orp��I�m�@�#�QOF���"�O�k����Oo��M{�$�]?��쐯2*j����)�8	/H�CȕR4,r�@��X"��BaD�8ZͦʧTwb��ɐ � ��
Lw���oC7(��<Z��j���'��$S�Nt��A��T�'h�w�:ճ���< :�F��M�:y�0�'E���N���'���r�$�ĀLC�i�Ek�%O��^(;�
=5^̹�7�@4[���f���Mõf��9�@X�Ŭ7X���S�y��9���d��#J����)�?J#�\hª
�C�
}��`y���O,��p�۳&H�$�O��D�����A��GKX����L	p9��ۧu� ʓ	����n�?�?����?)�'z7jE�'�?9W��1[7�dJ�g��J�珺b���8�M{2�i*�(�'Y��{�A����' �:�`G3@m.l��-B?�d\��M�
^vH(���<	0
ۜ�	&f�x�'�^��H�>;\H�<"9B�qǉ��G�����C#�����O����O�$�<!�b��b�H�9��Z��Y;���-��l��S�W�x���6���'�����O�`�'��i�FM��ӿ>{0�(��
�C�-Ta^m5-�����`�R�<i��φr���]�f����Z>����.�Ȕ�rbV�H�nHX��r�P���Fݶ?X�tr��'2�'c�4d�s���yǬ�3d�+�A�%���.����'�D�KdX�
�Oc�Co���dR#J�ʅn�$�; �)�8�cp��):�X�q�O���d���6=��HX5��)[��5O�\{���2�h\C!̓ )�Xk5�E�v-L(�'B����[�H+�vUnܱ��<�?����?��  @0]3a�^9(b�`�n/�?������||�yu��O2�$�O^����c,�J`� %ݚ�BKQ-�$ ���3�Ot!m��M+P�x?��%�pm�瓫��A��OB�hA���ݞ���s��N��|($ϋ-[����M�D9O"��%Ķ<A`�'[��A���R�\�Y��W�G^򫘒 |J9��'��O�B�'��R+�	���H���Ă�,�|1Ek�%�q�'�|6m�O�xS����O�to��w	�!3��M�G����m�9[�8b�4fd���󏅌g�n�c���<Q��-7 �֝6W+�4Bs1O.���O@{t�Qa!�X�q(Q@&�'�� p��!��O����O ��Q (}��'6�4�q��2@)����aǦR����WpT��?���B�<��֦������£�/g� ���K^Y���شY���ٻ�~®�3v��OU���TeV-ql]#pHߗ]�B�c�	P�~����"�y	#Y���I�nn��.O�����AA���x�A�6aPdMB�h�&=����	��t����ILy��0"�!r�'0b�'%*���a��I�M1a箕p��'n�O�}�'Xh7-��iC5����e�t��t��H�7������pY�U90O��Cc�F�~��|�Gˍ$^�2	��$��E��ͺS?P-R�,�w��" )X�?���?᳤,!洘�K~z��?	��%��)�/'�����oV}�*�:��Q��4�U����$�����	7D�Ӽ�GiM39�eHe�C�hbq�Mڡyb�ר�śCͥi,��T��4�X���'7䁓vo����$��.6� }s�aۅq�{ve��%D��;tf�<�u�'<�S�π�Z�2�'�b�O�ش9�鏵f��ip���UȊ ���Y��ɶ\`np`�ȟ4����p�8�ր�'ӄ)��\s�i�T��M��P�O�>���iu�6��H���OXf�+˟B%�a�)��L�V��7uVI�/��;Ϊ��!\�9���g����*B�)�Q����wJ8iz�hX�a��H��Xh��HVQ�@�
��?���?y����$	z� �Td�O�������@���ǇeH�q+��O�Pm�ן�b%�<?��U��i�4ݛ��G�C'z}�%b��u4��!��<Ŷ�w�-KN�	 �蔭�y�M5x>xm��w����|z�wt���gF*?ZJh
�A<k�戃'K�J{̀�S�'a��'X�D���G��y����[���5�8�q���y��'i���T��O��o�X@�q�4
C13@45"��^�$Ȃ���a�;�A����#�K��MϧZ\$�DL�J㾁�B�zd ���oZd�%��J�)�$JRm����XܪX�'�D�Dd�bE����O@��O�p���m�X�i�� p��de�O��ľ<)���()Z`ϓ�?�������3c>�Bs�s T!G��>�d�'��n�vl���7�X��D�p��Q�� �͋�a��T��pk@!ŏ#n�Sv'�f��Q��B7(�p%>O�D��?i+�>{�ɆS|��㝰Y	D ���ʒE��5��}x�� ����?���|:���?))O�A�t�  ]�Y��W6��r��(;�ry 䜟��ݴ�?Q�hQb~�(�>Q��iS<��a�I�q6��{�/]�<XE6Ms�Z1q�IX�Pf&=�q�T.���I���_w(��k��<y5k�>K��(�ēV�� �������r�a��Л�?����?��'O�li-�p�q���0P�HX�eX�<L�꓎^4[v�rv2O����O~�I�n��	7�M���hA U^x]�����>�\K�-���hڴ[�����'?���EDM�$(M{r����@T�i_��C+Y�w��"_��a�'���b�⟠"�.W��dVҟ�a�X:	"2��i):� еH���h�UxPl� ��Ob�d�O���<鷏�'b���͓�?!��iB(�k��Eب(Г	�3�fl���k�r��' ����d{��lR�LB���c���g�P���}3Ѓ�S�D�!�m�5�y�Ɂ�1c&o�F�ԥ�-��q�'k仲��Nk��2����dE<yGb����	���	1r��< $�]S�����ǟ���[|�Z���������DZ��ԠlZ�yǠ�e[���r�O��S�k��q2P��"d��8bQhB�[�>M	Ê��G�9n�FKtP2�R;$���+vkg�,�`kGN��.	�7k�h{�
�s�)#�6J�T�:�FC����8j"�/�4d�I֟����?y�"ҥY���P��*Wz@ԢV��=s�n�'��ʲj���y�'0��O rՈ�O�Q��Λ�$�&��Re����S}"�ȱlښ3�Ƒi�6� 8"��%�d��7J�(J�,�<^��J��t�Q����/@'���P&�03��O�� d��By2�O���Q�%j�' 
/�.P���9�z�hV��O��D�On��O�7�����a[�<��L<��4q�nD�v���IS�<���iH"������|}"bӠen��gd���^�@�F9�ʕ;G��	��
	0ݶu#��U;|��T���:��ƄrG�Sy��*��{PhǴm��٥�ѥ]����Hܕ8%
E�V���?i���?��'t���iO~λ{�P�c
4:��d���@���/O���àp}j����?YQ޴�?�G��<q K۲{�&����|@&W����+r��c 5�M�']������=E�z�ϓ,;u���?��rvF�4�$�t/�^��	�C$Ҁ�'c|���d�]i�M�O����OjAQr�	4drl��O�	*�����O��$�<Q�lS�A�Ը����?Y���
5�)�>!�,+P�hh�G-͘$�'��˓�?!ݴ�h���}H�a�
��?�i
[�^cLXJ���=ߊ�2�Q�Cr�Pq�8T�\U�p�Ь�VL�ژ".O���c��g�6IR$ۆI�!�ş��rH4o<��I��Sޟ���iy��9zBtP���H�Ɯ
������i�B�'О7M�O֨9����;.O�6�J����W� �B�N\	C KQ���n�P	����q����՟Dk�-�:��N܁k���'�,Qwɋ|��)&�P�,�(��
�&Va�x��'��'F�T�Y��S�GḔ
�@g"$0�wٺG(��,T�1������?Ms@�+Jv��y�,��3N�%j7H�,!,��c�&+�6���Z�������W*7��6���&]Ǫ��%�#�lS"��"�� ��)���yb�\�? ��K�$ճ(O���I�B@�Yk4$۟tk��%Rx�`� H.{�	����ៜ�Iޟ(��wy���$|y�'���'W�����;^A6|�&�ʵJ�
ؠY��B�1���XCyb�'���J	&����'n�*������~�"=;5OP&�x�5fߎ�yR�S#�$B��A?<}.)-���)R�'�<�Q�	�>%�r�+�̞�@]F�q��XN*��	�t�	��F@��^u�ş�	�� +cT�B�(�D���q)�]����ρ��qm�V�'���3�O�N�<a"�h � �(�B6dB�]����/Pm��@�
�3c>!x���6d~�x��@,2�nȖa�H�f/=�yd�$t�DC��0������5dԇFt�������	�?aQ�	7"Zֽ��	F�Ԕ@�,N�a�՗'h@UK�H� e��'���Oڔ��P^���U�̕@E)��I�r����T�[���$Fئ%ߴ����J��G8�L�ڌ��-A�-y��]E�:I�Θ[���Γt�4�z�-�O��W�__y$�O��.I��F�@����o��ȇd�#�� � M�Ob���O8�$�O˓�03� G�<�ŵ�	p��L7s=N�Pw��3"��I
�M��cӚ��'\�sכ�h�dy1e�+'�:T���A��9�f�P
A1b�4/�';Ƙ��<O��#[*�u穊����O�2��1S,�y��0�,����4�̭,(��r��?�?���?��'{�D:J~λyZ�q�/OP�:��p�"�%ϓ�?I�){��j T~"�Ө�DA�r�P}�9���ƽUd�Ɗ҉TZƩɦ�㟼��
Ժwɨ�lz>-���{����d�t��3ԅ�(����u/@�V���c��ҡ0A��!�'�j�C���<E�'~�y�n�����'����<J�.�X��W�j��	���C�r�'U��>n�ejb+H�\���D��.ǔ�`!�Z�%-��#�&|0$��
����$Q�Eyٴ�`���[�Fbj>e@����+�@;�HϫJ�R��R�Ǉ
�FJ�+3��Hj g~��i_�a���۴9�������#pe�=#��m��Ň�?�	��,��b���?�'�?)���$ٴ�2����M�4jP��kV$�&� ,1�ʓN��V�'D2<;�O~E�'�:6_4M�V����R�j�rq�>	��Toڋ�V� pk��$��t�e���O-Y��DX�P���'���aP��2pKV�1�fߡ��a9��y�2Ԝ	n�-ˤ�'���'�4�|��S,�$����9"�n�H򏞟q�v���� H����˟��I�?�h�C�yy�e}��-,�<���Ȍ�2���{h�3X7��n���M�C�n?٢&L1�'�Z%��$	(P8Y�"֐4PV �ýF\����D�<y3��K�(��ְI��e�'�&�d�-G$�b��O�pҰ��5;�|IsK���AJ���O����O.��<ᵏL7W?�����?�����eי(�B��ǀ%�P�)D����Ta!
 ?I�X�Tz�4Z�&��~&�U�? v�ɧ��E���j�N�G�te�$p��dO!-N�����\����S>�Z���O@�2�gH�{yޘY����S{N���!Ԓ��H���?���B*�Z@B����?���?q`��t"�w��\˼�C"��?I�@�E�<��-OXxnZ��K#�0?�;t.�A��,R�4k�B��cOf=@����B0jX"R�i�X("W�И5j^Fڞ�y��J�r���;��c��E�/]Z�&��?Ԕ��CD�/	���X
R-I�y�V�+��'>��'2��]�y�����VK�9�I�dh�SZ�0f��Θm������?�1�MFyR��"�2�h2�Y-d9�eӕ��w��y̛�}�:� @�O�u�������)�=m|�m��)Ƥz#t�:�0.P�}[����P�4�(Q;O�}Z�
��håc�[��I��?Ѳ`H�o��y���X�<X2��^�z,�4����?���?a��<ƴ�,O��H�&�w����u��$��#����L�c\�d�OV�DRj��O���?��4 Ҹ*t,E6��)[4��{Ҧl9����;b�ٱ �Ӵ�ع���f��3E�DI�
}�Eo��<Y^w���uJ&���%̳�f�@re�u�V��%O�	7v����O��$��\ c��&�9�)�$)ɨَ��G��8=Jܣ�I�<q��Z^�`�o�Tn�d��5��䊰Y mP�¦���� N�w���V�O�xڄ��B��6=�䠸aa����sf=O�쨗%]�(��ZpO�[yx�Q��+9_�a��'��l{�X�����
�h�Z��?����?sA­(E`�gMlӌ�J�����?a����H�2u ���OX���O��	�:{��i��#rS,�y$��{����в�O��n�$�MK�So?��\)p���!��{Veי2���o'Q�������vuz���B[#��O޺�	��2&6�S�\����a_�uuj��J(Ht�Q`QgB���J1��3$�Oj�4���d�Od�?6N��Q"�}Җ�qҩЏ~3�E��$1N�z����?���i:r%H5����Ly�ijt��W�\�����q��4P��
�fw�l��&�Ӌ9 �f�� o��d<bFi]w���+�C\�<A �'J��2��[�V��|�c�S럄���&��c��Ц�?a���?��MKt��ʟLP��̩z�-�K��<�`���MA�L��'���'���#���Φ�]4��0"�N�@��H�˫N�2T`۴B��g�%��A�`W2�Q̟,�*b�'R������f�+e[�Et�-H$�1b��.<�69�EU�AS�S�D��1��C�G[�?Q����p*:9R6�L��ꨘ�iV�?q��?I3DQ5��D�?�����J���Ox�:��P�\&Lq�J�0fH���On�*�7O���<���iD�6�ˎ�~Ll��u춤�� S3, !1%)C%��aW�S� ���Iuo0�g`^$q��� �{���;s��)�I\�>x���C53��hY�����
��S�"7r��'�"
E�l�E@D�'��g>k��Ꮋ;9��u�L���R<�`�ai1�2��2_"r(��O�Dy&��O�ؐ�0O�	o���!�iA�W�ܠ�֏5C��!H��&M)���'bY�M�G�X4_4�e�W��+6�~�B�k�t@s�=z�H �G�EL1eH�"���چ���VƔ�'����ݢc_\ ��O"���O�����u7�8�M�;k₹)���.��$H&�<i$U:bWB�e�F��?����G���<���R����G'�1r<�! ��"�p�O��h�FR�ϕ��D$z � ��?�h��, �EF�DE�l`�M��d�P�H1@\�]�H�I�3,h�i�� �D����<Y��'�f� �%�2��i܍ȤA�!K��A�Xd�w�'�r��a�R`�9 �R�'���Rㅐ$����wĸ�jV��nY�F���ybc�\��Y�yҫs���D�O�(o-�M��)"/,$=qb��?}˺Ų�C��t��sUL�"�ݳ%�[�?a&�8)<=�5"X?o߲TΓ�u�K����C�?�ؤ04F�' jXC �K�w����`̕�?����?i���dȡM~λQ�
@�3� �	��� )��D�S@߻�?I��=C"�#eo�<����?���X�Γ@�|y8Dc\ Ox��!cI�/XN�P�kȼC5�F

 �z�ҁ�k�Z�I��'�&��,N?MK����!�I�2. ��7��na�3�5+����/Dp�	�?!�/�@�*D���?I�O��ȉ�5	T!��MMs��x��?a��
&*�b���TM������?���
zR�yQ	D5�.�˓�����7M�#�����ĝ�@��?1G�i�N7��a2h��*݌�������.�r�o�!�X�a�ڤ t}Jv��C��z�%��dv��0�g�OX��N{yb��s�Щ07g���������'d�BS�I�������'��\��{�dͣ\�y���k0XŠS����cF(�����	ПP�C�3�)O��mZ�JZ��B��8W��㐏\�2j�%��41SPo�DJZď���?9���et��9���"ڂ��+⬱���+���n�9=���	%�?���69��l�<�'9�n��'ǎ$!f�i�p9��^�g����h�$y�6i	]���	�?��@.�T��yw�(,0�a�y��d�rL�4Y�zU8��i�86��\���k���ϟ)�J�^�8����~p���
�ͤ���ӏZ���ѥ'��4��N��}R�T��A�S����L	c?q����O�\���ɔz���`�"O4��1�R%	�ʓ�?��ҷ'ͨ�Q�=�D�����?q��}~"��>q��iʦ6-��N��d4/T���`Z�Fs��&I��6�N�CbZ��yB�H+i">7��	q�`$���'?<��ɹ&{��+�C��8�ÐN8h{@�;�G΂��'b��,�0<P�Xn�.ce�o��*�H*�?�$�Cg�
Y����?	ѷi�bB� ��4���
q韌A�pPFG�w b��"�����:A�ɦ��weֲ^��B�E=2�	�f�0q��k,J(?'ЁjC��	KY.�q#N��6E<�"��<A��'��R��ƍ������(S|��sf�Bp�X"�xb0:�O��e��;sD�ʓ�?Y��/�X$�O��B���ԅa%I_8%����l�>A��i��7Mн*���R�n�v0�ȟ4���k��Wvl�g	���ES�mU��0�S�F��}���3S$l���W��aA�W�l��r�\iB�?KLEC��^�k�
؉�$F�&$H|��ɦz� �@dMҟ�Bco�� ƅy�*�xF�e*��꟔�ٴ�?A��a~r�<I���MC�f`�? .@KEy��Q�AêD�踑�l�Uh�PB����$�p�Dk]w�q��nP�c���D���$�!8b[ jwH� %��|zm���4�zi�B�ɺ��bQ�ڗ 2�A���'V�X�|t�zϟ�lΟh�Cf���p�ތ(�,tq�c�&Eҝ���E���	f}L=����Ŧ�S'nX {��ѭ0��I�8��]��Hr�8��劇1� �@#[x�+ԊE���}�R)�*,Y97�'B�'�u�$�4=Y�uҥo^�F����'�RT�0z`�w�l���П��I�?e2���.Atqig �u��la`ƚ'O�����I�|mڗw����	D��`bB5����ׇXqN�Y�rMذB�ݯM|@�*#%F'��28O�$HG��?YR�y��I)�1��,kR��k��Z!i>ey��9�h�X7d���?Y��|r��?�+O<�"�8d<Ttّ��q֚<�A�v�l3�<1s�i��$R�����s}�r����dk��?�|�x$�0->�H23 Ϧ���} d��/�) -z��-~G8�p���2�+V��y�9D�� ���-��ݫ����?���'�@hb5��<���'���O��A�_>�����&�l5����<< ��^j5���-�ӟ�������(4�SΟp`���;���X�h��^;`D4�����)�JkӬ	�U�O*�O\���i�h\ #�GI�D(`Hi'(F�N�")�A��*{�
ͺ43Ol��'gѢ�?�G�Y%#�I��?�'@΅gJ�X���+��	fjI��4CE�o�P����?���?�,ON)z&HߤM|�D�O4����.��%P�0p嚝r�D���O�;O��$�[}��x�,�l�7:�l�		b$!d!ו�� p�� O_��1�@�v	�3aJ���ƞ�L��C�_>�B��O�:�"��k+:9������� 'O�
]hL���?y��r.�!B��'�?��Ӽk[� 8��?Q���������	�L
����ڟ$���M#����-��?�;O؎��f�V�D��S*v ����Au��`C�i���7�S:�Y&��9�y���y�|�;lB�z�P�/��RT�@�)��,+-�8i��}e2�F"�ZM��'���'����9w�z��[*^@�gCB!ka� pX�X�bM>F��I������?�u�r>-��j�,u�FF�,���cN�&���Oram���M���V?I4�!pK��e �*��ŪD���@�����H�iI�	�ӈ���y26cE�l�Ɂx��2*Or�	�-F4$@�*��NI�i��(�5W�d� �JK�U t��	ǟ��	ٟ$��iy"K� aRq���'X�A�cQ�F� �iS�#r�$%�%�'l 7��O���E1O���b}§tӢLn�r�|�Gd �1tr���p� �a(	?�:`q&���4d��I4�d�'��]Q$�������륮�^q��R�IA�Bf4]"Sc�NU��L�L�����'X�'?�� �4:e�C`%����l�!�����	7f}�B�s>���M��t�d�X~����(��@�!�J���Bn�o��d˶C;����|��)�E��So�:���w��B�%�M/�U�f�(*&��A%.�y�,�\��ɪ�?yf-�Lf���?��'Ǽ)�V��N�ڡCFgJ�}���b��?�.Onm��I]A����O������!�5�M�>L�z0�fl�dq�	���d��ٴ9��A�$�'���6"�|�֨ˑXy:�����0H"Qx�O@/kB@��ێm�����<�./_h���%>��D�'G֐B���sݴ�{&�	�Y�����O��Q&�%�v���O��O���<9�hV�/ݐp��̂1�p��̗N��X"eR~�}�8���:S���6���	��Z�
.d�z����R�u�`�j�M����1�J��d#C����]1�#s�z���q).�����hY��b�+�� 9�g�!5�A�O~U��I�����O������d�|�ቡu��Qx��y��!60(�+���<���?!�'@=��'�"6=�bMH ��s�r8��cͶWC�t�s%�Ŧq#�4L�X��'x�����s�T��5ݸ���n ��|��c��
'rhݛ���R��k�'�Y�%���� ��.���	͟@S#����҉�I ���*�cș:8B�nˎ)���柌�	���'��Z�Hݼ�y��'�R`�0'V!"U.�= -`���rB)���D
p}B�aӊ�o�	YؾI	�`w&˄e;H@�P�^*)����È�|���Iq(D�W�Nd�a��|JP�ʟ��'��9;�4 �@4)x�I�N�@ޘ(4�'K�'�z��`^�d�O����yǠЩ�'� 
����MU,q҅X /����O\4n֟,[��=?�;I��| �-�N���A"�0G2�@��a$h���뀼iC 㦅�q04���/R�y���n�n��MP��z�L��RK�ْ� $E�\����[�ܘ���P6>eT���K�d��ek�[�}T�C��1Q�9��^���u�ч�|� :� ʖVOL=�Z� �@[���Eex<ɵE�a7�իB�̸\9J+��Ir4�!'����M/I`
l�Rɜ-h*�-�ЩR�KD�Mʳ&��*�����'��X\�j󧄎<��M��@�(�z��ݪ Sb ���Q���u�SA�F}��N�q�S���j�5�$���2b	��x�`mI �T�g��r��N�`�����G�4��%�IF�X���Y0M�4��\����,]�<�4� -VЛ�'��'��De�<����d�X}@D�#0���a�$9?�>���ǟ0�S}�t�'ɧ�	��N۰a��d[�[���dA!˛�ۄ@z��'��'���V�Z��x>-��p���膢Fq V���4�?a���1ה#<�|:�,E�',X�f�|�s�
V	'�lAjf�i���'��dJ�g�"�'̶���O)�L�M��L�=8P���`d�����'˘�A3���M|���?	��E��u�7�
�tٲ �3*�@82��i��@�mIR�'b��0�Ok���~�'x�8�qfĖ�@!(*6�ЩE��X��x����$�O��D�O�D�O�A��5g��a�3jZ>,Il٫G�׉�4˓kb܌���?Q��CB?�S�|�k�B��(�o2���"���j���ٴo��8�'Y�'�R�'��oD�0��)�9#��ԃ��%v��SF쀸G�&��1���'�2������y�'8�`l��D,[�f��J��c#$\!"^���?���?����?ـ�����I�O�� �j��E�a��ق�	�; Ӣ8���i2�Y��~-��?i��z�RD�	" ��@�
�� Ńwڳ#L�7M�O2��<	�OO (y�O&��O���� l��{Rt����M��mBJD2�~�M�?��P��3ʓ\��0QQ��z>`��ǀj�\n�Vy��RL� 6��O��$�O^�I�@}���1UTP����t��E0%gߜi\Fl+F�'�bm�O�a���x2H�6���I?y�8���2�M{Q$�3A���'���'���J�>y�f��<1���7Ffd����K��!��L����fΙ{�r�|�H>�OI9Z�����$��[�8�[&j�_1�6��O��$�O,��(�]}�d\��yZ�M�$ͦ���ń){�j����2�21+6B.�	>&�2c�����4��rRɪǢH�CD�B�J�N�P�ڴ�?!d�ιL[�I�
���I����Q좟���Z����Ϡ�&�ݶ=B��1R�x��$Cp�����	���'y�Q� 愖.�����+�U�Tp C�6-�H�]�*M��?ID�K?�S���I�Y7��{���6_��E�倢
`Œu��~��h���h�'W>�c�%v>�rPmL/!"Y��Y�w����$dnӠy�E>O �Đ<U��$��@�$�OL�Cd�h>��"¬
1<lR2 �%�4�hGW}��'D��':��"X�{��|��,F=v�2U�̥!����5���`��0m�ΟC��D:�E�Ov��L[���0�ԧт�d���Kv�A���gӖ���O�˓{�����X?�����S�F�:�K�bW-UR�����.CA�p�3��� q�
�Ov�Dɾ2|��|2�w�8:U�M�R(JXQ�ߊd]����4��SEG�)oԟ �	ϟ������Ф/����+�v
�jtX-6�]���O@�d�i1�� � !�BG��Ʌh�	j�(*Wg	�/���%+}7��O����Oh��b}B.?�yR�H=�-AGn�`��'h�Q�J7�/���Hb�:��쟘I2G^�v���eÊ{1<� ��U��M���?Q�n^��j�Y��a�'k�t��k6��2l�M��f����ي��OrT�� �d�O���O����ϙ)���&�>H80�������I�9�F�ʯOR�p�>O����!s���56�p�t-�c�
�y_�l�sNC�����8t�O@�d�OH�D�<�Sj��9�9x`d�'4a�ЂWT� �%^�Th��`���	�}3d��Z���O�}(��.L\�
0a�6r�@�!�����<����?A�����\	���'{����D�k� ��iF�Q��	����Op�7�O��S��'�z�hge�;��HTn��B��Q�L��?����?�-O� �Х@�ӕ�L5�Jg0{����p���ܴ�?�q�BE?�0�My�O�����	1B]IE.�eI�D�-P��?����?Q.O�A{㍍D�S��$��'�ָ�F*D
O8$ٵ�L$�N�`v�O4��P���_wE���9O��z5RXd@;D�F<zv@�������Ȏ������� �	�?ݗ'��p�J�{u�}�A�W:t{��Y7d�B7O��8tN��O�Ov4��fH�1sN9cjM�İ|�ݴ�6U��?����?�����,Q9�϶+�8�iG듵|C��W��G�<���#$���0��)�'%��bpJ����s�B D�)g�i<��'m�Ȓi��	� 8���<���z��Q'ᐪ|�D��"��_>��a���g�'3�c?��I@?��Ͻs�4��RM�v$m�©�����p����'��$k�O+�D� �~�'>�\�1����Wr�;A��*mzQ�p�x�m������Oh�D�O���`8��4�|��3-��Xf̓ �/+(�ɥ|�
�D�O��Sמ?��u7b$��D\�eb��i$�M�����d�ON���OT�gW(�s7�Ĝ��B�74�`���[�d�8�'�ҡR��?�5`�v?��Zy�O�����Q�*	��D�%������!͎��?����?a.O)��LP��J��Q�g��8�E�Ag�/y��޴�?	�kB7�yB(�
�?�,���D�O�	-��ŸJ\/m-�3rhC�pq���'��]�|�����ħ�?���d\W$4�J3&8h��ЭH-/.�D��H���#h���O@��?�i݅���5���R�ׇ|�r]��F�>9����\����?9���?����� �2��a����xȇ�
���OT�I�S��e��)�pKb�QQjʱ,�b��P�lM�6�Ѐ�L7M�O���OB��BiybD�|
���M�*|�GȗN~H�+�%S�q囆��A�b�'Dɧ�9O���ۙBL�9�ӨB��8z��r@��l���t�	џ,H�d�
�����&j�D�Opl�'�i�h����B�U|�H��&XԬڴ�?9,O�%�5O�ß��IƟ����@&����t�B�Xw��M��?F~<p�^�`y�kv�|�Ic��I�?�آ ~H��#ƚ]A�*Z�F*F�*������ğ��IkyB�B����FX|�r�"L&�&QQ��>� \�<1��,���R���?Q��(-��7�ʘA,�Ḃ�Ǭ;���<i��?I����/&�>I�'�(�!�n�# �CIJ<nڧj7��ڟ<0��y�x�П��I-n���C�$@"b�<nN6�[%��Dn�ԟ�	���Qy� �js�맧?�� \o���C"�v�����_7:,���'l�H�'�v��W�'�a�!��4���FZ42~@��A�1d&�q�5�V��M;���?1.O��J�)�Y���'��O���@�蝿}4��
W64�PASR�
�y�gNw�R�'�`�'�Z����w�Z(��:?�V��ũ߰c�:��4��DY;5��oZ�� �I�������� f�? �lJ^!(��=����lG��[�.�	�?��XL̓�?Q*Ob��������r>d��wHO��$@Rc�8�M��o��L����'2�'V��>I@L��<�A�Z�5��J�I�4�Q��%ϗ��6-H�y�|��_���O���/_����GZ�����v�7-�O����O����q}���y��'�۴`T��G(F���),soV��Q~b�)r���?	��-F~�)�iL�w!�mI0)1l�&xCc�iR��#L� �0�M��?W�E�<	���׃�K�Z��jϸ��8z��e}"���y��'�R�'���'|�I�iW6���m��&R|qɖ��C�x�ӆΑ����>����O����7O����O|�ܴ)��i�X��8��Y� L#�5O˓�?����`S%pr<�(1��&�/y��A�@��^����5�i��'x�JV�y2�O���'�q�O<�z �́%�\��K�prB�_�Mk���?q��?�(O�Ѓ`�D���' ݑ��$u�U�TePѱ��s�v��L�s��LJ���D�O���皟���?'��z��4_1�J��	A�i���'�剗@�M����$�O��i��<1���D�� ���#N�QlD)8T5OL|�q#�O���H&���<���P�Q����D҆>�*�󧥔�8��6Z�k�쑐�M#���?���ҥU��J"@U�N5��T��eP2���zo6��	�,
�q����Hy��	��'g����'�Ç=,�a� �N�z]o�?�l���4�?q��?��'/���|Eb��=u� <)G�'5�0	�p�ص"� ۴,pΓ�?�.O���i�O2���k�<X�WV5>	¬�"#A�']�&�'���'����u˫>A��<��R2
�n��atBaѫǈ1d��pFC���is�[��K�e��?���?�J�:����U7S���"�#D<p�6�'�v�(ᅷ>!1���<���&|�pϓ��1.M��ek�:�Hp!��B���'���'��ٟ���ܟ�'2,k���F��3	�>h�B��*rZ�M@8͓�?	î��<��'�?���g!�R�'U#GᎼ���)dNl!U)�w��?���?y��?�熚/&�������SF��$��X8A ����6C�K����O(� ���O��9O,��b3�i�R���[���[|��9� �i�����O�$�O��D,I�]?-��]��P�ɀ*18��6���#��iڴ�?�E�P�<�DP��?!��Y�����29Gt\�U* �;�\�Q3H�iu��lݟx��Ky�%�%�(�'�?	���RqiIa��!��98d��Սל�da���ш��?�E�SZ~2W� P�w�<���^+d���Kŵlh���޴��$[�f��ho�	ğ������M8c>�Y�D��/wG�Aa +�;v*^�;W��O��d0����O�)�O�����(�:c��P�0%H2k�R	3����MS��#�F�'���'��D-�>���<�f��%R�>���2I���Ӈ˄����%�y2�'}�ɩ��c>I�I��Q�&l�/S�"A�R�4�
- E�i�r�'\� �!X.�*b��$��Ej��s30ZI�UJWX�i�$�3�ih�'��y�f6��O���O�L����M]���`+��]f6�"�FFߦ��	*H}�j.OXi;�'���S�����r ـ��oEj��V�isl�P�J�>q�e��<�)O<���O����<Y5���x@�[�Dٷ:��`Q(��2��dJ0T� �+�O�h�ʟ�	.Pb<ȑW�XBJ)j�&��5��P�e�,�'���'F�X�DB'�����O+.��1��m�����a��?��^⟔�IF¶�	�?!�	ɟ$@BE�?q��"v���%?���w�
xO���?	���?q*O:Y����]�,`j�pY�С	s�G0@�d�X�4�?� kGM?��ECΟ��I9;�����q�D��'@D�����3@k@Z"ʛf�'��P��q�E�)��'�?���/�!�,�9��0 \r���#�FF?�rɍ����IY��"<�35�.�Sh !B*R��	�
y�E$�ia創o;���4V����������Ϋ5��)���`s �KN�p�'�2$݁
�O�2p����۫Lބ��DOtt�!+��M��e\�&��v�'jb�'��T+�<��}��z�JP�T���k^2@Hj@�2!ބ�M����?yN>���F�'�?��`
5l�$��3�|�$+��,iS�V�'��'-Bz��<#d�0��yW�7�ԫV���`��#}h��Ą��U2���|�!š�yʟ����O8���72�i���C�0A c�
�$�oƟ �0Dӧ��$�.�y��'�~��Οkl��dݬ��i$8<4`� D���I�:� ��Ijy��'���'��8 ;u���D=@���r:�<r�@\	�� -���'4���͟���O�� �ЬCָ�����(�	6Ȗ-:���<����?����D�7M���ΧH,T�QB�jxp�`���k=8`�ɬ	I��$�O�є:O.���O���W�:�S�����@�x	�0��F'T��9�'�"�'`�]��9�]��ħr���03��*c}"���B�R�Zsb�ir-�~"�V��?1���̓��9r�<[�"''��U.?R6��O��Ĥ<��NMP�Ok��Ob��q���#�b���/�%}?4ͣfk���~��8�?���fՖ`���[�n��x�pbwc��l@�#G��'Jכ_�Hp�4�l������O|��MyX��ry��$Z�rb�1+��vԬq���?)L��<iO>!g�w��(5�dZ��Y� ���y��=ʖ7�Η=F4o���h���X��6��D��yr+�7)�F� 3iM��bx��@�<Tf7m�A$��9�����OS2�
��&�	� 6�
�.o��6��O��$�O�1ZRk�Py&��<��!�z�o:� ��'r���[T
Y� N��гi|�' �S�����O,�d�O�ġ1�Z
FV-����(NMfq	 (̦U�I�^��u-O�@�Ox�$�\��i�H 96��Ӯ-���ӗ-Ʀ|kI<i����O����O6�Q'���� ��hɴDj��C�Vu�dhw��K� iX��u�3��?�Ik�H�/P�|	���9.R]��N�ͦ�����������؟ؗ'R�h"�f>�xC�V�&l��� !)�������O�\���'H�ă"�~��<I*����ޭ&e�D"iC#����ǌ�[Q�l�'-"�'4"U��q����ħ0�z<��#M%L5r��R�!�8���i��d2�~b��<�.�6�#}�	<&:���4�Lp�KE�I�M{���?I*O�y���S��'��O���A��I?��6
۫]�È �y�I�&��ܦ��b���	hy��c�=��b�$*Y��x���!j0��q��XʓlSf���i;B�'Xr�OG0�Pz,86��"2�:CːA���$O�=�?)�Ta�$Γ��2P�l&>)�Rhک8�Nax�䓙7�ad�oӴ]�n
�E�Iß����?�:�O�*U6O|M3 �^� ����v��F6�``�ܦ���e+?�(O�MR��)�O�M����7�PJ�I� ��5R��Ҧe����,��(e{ �[�O ʱ4O���ܼd��'ʶUm (���PJ�A���'ҒA{�y��'���'�V����,z���sE��|Qv%A��zӀ�D$D�^��'�R��'S�KG �yr��5f�J6�R�afBܚ&���c���)�M;�dPAΓ�?1���?���?�/O@ hW�_ '08)�%Hrm޵�`�2+�
�'JnM��'>b�T��y��O���'�x('f@6)��"����2�"�̕'�2�'}�_��P1$�5����� �¥
3A�ikF!�Q
2�M[��K�<Y��M�v`��B��?��Y}��F��̠��a�[���B�$��M����?	�����O��"A�|j�'&$�Z��(!c�D
dK!i�08ݴ�?��L^?���Fßh��?��7��C�&D�3O�p
U�\;Ĺi���')�əhR��O|B���4o^�Y�<a� �GS����/W1A2��!z�=���<�,�Q�|�$��d��+\$ҩk�p������륾i� ��?���"���B �`��r��ػ�MǁM��$���Ob�3Ka{2k�-#�&q�cK=\��ܺ�ڂ�M[@� �v�v�'���'��T��<�AŃ(2� %��	����f�p(���M�bDT�'� ]�y��'� ���D�<w����)Q��3�g�R���O(�d_�fL��'�`d���?�a��æ� �� >U�Xj�i֨%�Z̰��2���+�6b����ɟ���O����@�Ղ1�x�j�O����ܴ�?����tq�OD@��;O��ĉ�J��d�k \��Q��,Ű����	"'���?���?�������lA�)����z�R�*EM�S� A�u�CR}"*_2�y�'p	�'����'���I�#�@%!p탧/٢A�a?��xj�y��'���'��	�(h��p�Oz��C��>.�$���*y�X ۴w״��?�E(��<q�'�?I�JCz��'&�)�%@?��Pȵ

!	����/O H{���#�fT�B�	��~e�d��C�Ɇ>�>�[	Ե9�>9�q_�z���	H��ݩ�)	?��s��Be�� dؚt���PcNK5aDpd��k��E2��gD�!�fl	-]����\?=���#-Q�n s���W�����S,���j;q�P��4�%2�[1�Tr;���@�=v�* �`� oX�������<�T��7X�2���f����O�ٚFDjػt#R�pn��"a���M���#����U��2$�ve�韰�`s�(M��� �BTQ.�9QN�.w����f�N�qhdY8"Ŵ}{�԰�?E��n�Z�� �66�B홅�I+���^w�p���O�S�l�	*�z�B6�57ؖ� &n�1a"OF��"�Z�/
Q�P��4i3�m�6�x�G|� !* ��?��[�����ô9��\�4gF4W������?����5Lz<A���?��?�qK��Wߤr�Veb�;�)�f*�ȓ/F@��x�g��*2Ä�O�����'�p�*�	�&K�e{��68����'��{��փ����b2O�yr��e�:�`! [,"P�b4�O"$��'���Fy"oO�|�P)���7,#���a�ρ˰?��>OJD�d�^�I��b��ڑ�J�k�H��>���	z�T�'}��(�9��Eq��Z� n^�S3)ɜ�P�!c��O �$�O���Y����Ф�O��8�n ��%�Wո�!�"ٵ��X�G�;Q~�(c����=Ɇ��5(lI�SΌ&?ܹy�kY$A�$��h�"=�����'�5c���?I����|A2ܻ�N�55���Tlƛ�hOv�?1u��!^N<j�(��D��9s'A�~�'�#~b���!{�P�2f�S�r�\��1FJ�<I ���<�}��5s�Hm!dl|r�3X��(!"O��cPMٚښ9)�)�)o�4��"Orx���vdt����CՐ	�!"O��C�Z��$*`��t�1��'D�t�m�A�;A/OB:�I��	3D���1$�<#\4x�� T*V�{�/2D�� ̰g��aC��9*�:)�"O�#��	�	������19�"O�|� �]�g���ȆS��"O�${u�.̬D��@E���"O���-phU �����=��"Otq  -І^B��0r߄E�e"O�!����H��a q����S"O�%g��?7N䵳v!���e�"O&Y��	M�s��k��;\�q�"O�u���g�6�ɡE�КЀ�"ODu�3oG����1D�v'$e�"ON�B�՝<�lp��X	U%d�"O�eF�Z�h����LB��"O %Ш@�G�Di
d�Z)X�"O����C 5 Ѽi�s�
N9�Y��"O���#q b�c@��2#��@�"O"�n� N榄���x�0;�"Ox[C-��ϔ�K&�¦:L��s"O�໢I�f:�M��n_�6<l �"O�p�6h#C}��ԍ�7���b"O��)v�ǆx���	ĬG��4i"O�� �E��&)�p�O�v���@"O�Z��ϑ|�$�&�<,���"O^(j6�N�'t0 ��i
>@Qԩ9�"O����6Y���<k$js��yG������s��e��l�B�H��yb��������m
��0�)5�\�y�
�!#�0% ����u�
U�y�DQ��\=��"�+U�T��4f��y��RB9����L�|��c����y���C\Й�;F2Piض���y��:OT�TAʒ�4D�;��i��5�F��d�	5,�ޥ0��V�dl؆�s[��u�T�HR(�Q!~B��~y��T�W�)�B�ס� e�Z`��5���a�����E���߶�Ȅȓj��
���۲��ѥ�z\Ѕ��J;��49���#��/l`P�"O���Pgݐw��)��B@�MFy��"O�]X��O��Qt+�nґ�e"O��Y�K���*�P�+Qp�2)s�"O�d�@"�-�����W�jMRɋ��'Y�	-OƭR��$oj��Bl�6��1��"Oڥ�282����j[7g���3�I�8[
!F�Ԣ��d�	s���CK��y��ذM���q@K'���r*Ģ#Ȟ-���=�)��4A��c�Z�:��L�Af���R�2D��,��}��%@�'I�8�<�cb��̳, HX��k�ŞM沙i�ꅻÀ$��	0�O,CH�>�� �V8�S�
�����b�<q��K�G��)�F�:RCs�T]�'\�15�S�u1R���0┅8�l�!-Z�B䉡( �I�f�(b�j� RÃ8�6�4��"~n'��t�L0�j�6��LQ@B�	���ѧN
0�h�!�[��C�I>9+"5b�C "Z����!�?��C�1A�Aw��?��Y�Iċ<`�C�ɂ)}$%��UPC�Q�#�!Ԋ��$֋L���<�"ЌJ~Y��a^ep&�J�
5D�L8����0�(�Ja�ݞr��h(��>��R�}�Z�b?�xw�V)h|�C�/LQr]IЁ1D�`�bG75!��W�U�m�pa#�0�I�-pc'�'鬀�v?Txڴύ�*��z�'i���Rě"�n���K0A�H�Q�A�+ż�#��� ��'*��<-�08DH@�iP4���'��k�����'��]��g� s�0x�;z�\���'֐݈R� +O}x�Bp�ӥ\%��H�O���̇91O>� Ǝ�)P���j�KD0%l89��+D�Lz6��~���� ��9YS�ͦc�'�:�q���y�g��#n��<ja��PX�3ǄA%4*�C�	6_�X��O�Zn�Q3��)VAh�bwM]�a��~M�s̎t!���+��k&L �p=1u�'kw������84m���1 ���7~���0`ӮS����:��@���:�XhC��Z��<G
�[JȨwD�h���ǂ�֦���&���ꉨ���#�-�'L�`��"Ot!:"kT�P���c+�-"���5A�g2F�
�(X/~62ܠ%�i�6#|�烈D���:˦p��KӶjm�`�&%D����*X�~��B!����O��a�W(�4�U�ȡN����I�x�JXr���y/:�B��X����'#Q���w��* ��� �Y�8VJYp��
�9�:�@��H�E:�d���Y�H�0�U=J�$�V%W`�уT-^�~r
�J � ��0Ax�R �a�@1���nިC���Az0�Xr����0�Z�w��* �p�޸�w��	k��m��S�&��F`V<8�W��.JЩ� �~�D���9��'��@���y}��v��J �$租@�����9�.��w�KNB���.&�l�´�G�_������H*>��Ă�%]�d�d)sŇ�77^����Ɲ	�������xq��K�19lݛ�A۬$id�>1Ea��!��PňU Z�	r�G�<Y�̐1Y�X��T�$l�2Ai��aB�R͘7�Z�v�W�<���D�M�j�*��E��I(�E�[�Lu��,=�O�5���"@'n�'++Q�!�Y!OeN	S\���Q�낷Q8�RW������8�P�w���RA
�O�>���(6@��)्�>@��#DC�5���%�%\n��M�dq'�� T	�r�x���֒����C�>1E�?����i�(	����I�P�'����Ǡ�9<K*�[��9z^"f�^>��)ѳ�9`�x��ҁj@���*�2}�<���G/(�̑*+џ��g�E%�Tt���u���3�`��ROD%:���	/;��c�U,e}Tu���5i���7�p�xQ���l���P��$(7J�`-�7����	�6�\���_;$����3肔Lӂ�+� ϕz8��fcZ�}>i��%	�v��O}�i[�@�W8C�"{�蝌?� �{P)_l���/��}+��20��9S��� >��m�mĕ&�A�.�$ʨk�F �<'jv������ɱ�l�c +_�i�DP �N6��">y6"��}p�k�͝
n����
�#�b�
��HJ�3׮�"c0��qs���� � �T3m�-0��=w'8X	�3�gM�,z��E+wպT �eI�"�J͓SaJ�2׭J$R�i2�E'��-x��U7U�U�mY�bJϓV��P)�ӒP��,0�PA0-j1B�b_0���2��xÙ�'�ِtdy���a��߬���9�Ɓ/�V���<r��'OV��8��|+�X+�h
1�?WפQCP�'ڸh��Z�(����U��!sux�q�lK!_�(cSɪ�9pS�x®���q�/t�l�'��2�~��[��%1 o+q��ܨ���ĈO����߾ �"��Q���ӱ���pB�n��[�
�|)<�D.g��p���X�5(`��ӑL\Q����L���e��wB%���3LO�찂E�D!�|I�aHm�D�c�`N��j1�A�~���(7K�6��p��m[��:�lN0��RÂY"k�Hd�<QǊI+0Heв�K�O�e�b̟�O߀�X0�O�j�P�IK��`]��'צ�p���s��Ԫ�K�'(5Ppe�,G͎�:�@[�:N��t�R#�(�(�P�.�ВAT(k�P)�*|�D'�$A�)�(��$��T6�d�}�H޸�8�ig�(F�\�0�J��<9��C�6���`��U-.���dǘt3�=:�� =U��Kb
M�W�f��'�D�R4.�+0�N��|�&�pN��5.�,S�,�@ ��]���&)��r��U2�2���%�2E>l	)�)Ϲo��g�9)Y�dS��Z����d�eK'D�-�Ji��'��}��$��@���&6Ɲqs�_>T�e�牅">ֽ1�]�P���B�|L�L:}�խH� �>���Б!@�q�Ŭ×�~��H��y�<)�>�w�F�O�X}Z/V ��K�H]�/7?���O��%A��#=@�݂XE�X�Of��8���#��,�QؠE~�x��H*z�x�����0��ɐ"���E��hQ`K@ȨJdiSdCP�f�R�鐯5�~}0�a؝Z�<�.E�Ny!��Y����"�@�m~\a�/�5j�k�m�d,V�i�*��I��UMEx�NYy7lF�#��`F�Rt�<���+��J#��^Xα����h���F�N�t2�O?�DD1��C@�),��(x�)d�!���a�V��Q�� j4���"�ˉ:<�	�Th}�����*��R�N>��	@@P3�`B�)� �ܓdKW�o�A�c��r����"OЍ���)xl,X#͌�"f��"O�xy���5;�A�t%S�a[�3�"OX 
E�̰	��h�t�Ԧz� A�"O�EI��$l��,q�j��/�����"Oδ��,n�v-Af��9#��=�U"O��C�1`V��pgN�L�� ��"O<�"CQ}�v0���~�R��"O�i6�_��z!Q�'�:z Q��"O~�SP��V�kSlY�QR|{"O��sj�r���(���zU\��S"O�m*�B��z�l��mH�NA����"O�e[�B��T
t�C15AB=�"O�1I��4U�CNʰx7�u��"O����kĆ[��{�OA3 -6y�"O���4�ǄJ��I�M�*�h*�"O�WÊ;Z���&l�E��ͪQ"O���O	$(E���\b���4"O�b��8��ϝ� ���HR�<��)�!h�tA��(7@��R��H�<�"��� ��C��31(���AE�<�vOY1sN.q�nK�&�(��G��C�<I#��eQ�1���ɳ@��$��RC�<q"�܋s�́y@�0k��3 U}�<� �o��°,����p�#�x�<1k��hO(�዆:-���BBr�<	&O_7���4	϶ �$�JC	�x�<�蘫6�@�ٯ�D)b�$t�<�a��u���IC�JYK�-jqˋo�<����]@�J�AU
뎴�S�v�<i�O~�hS��)?�|-��/�g�<9�F-��AT�ɼ
]Ա*���N�<!B*�kP�XDI�dv ZT͆I�<�+!t��	T,�lf�J�J�<��Дp��ȑhR���A��~�<ك�c`$�!]�>�)Yq�z�<�q�����$�R퐱9�nI��v�<qC-	�b[������0��8:Ʀ�K�<y!���\�����Y�t�i0I�<��o
�� ��^�Z�xA���F�<��f� l���
�.y8 ���@�<)�!�6K2�\�G�X�Y���pvfA�<�an|�F	A���!.�9 �kJy�<���F�NȠE���-�0xQ⣁m�<�UL��,���`PЎ�p���k�<ق�߁/� }���]
-Q��g�<y��ΏQP��S���<��f#^Y�<	�"f=8�yD!wwN��QX�<�`��3oͺ�Q�˜E�����QT�<�5�Q9G��A�uC�)���xp`�O�<��6 �L�Fe�T%���l�O�<�C��'#6$�i����L(����Bp�<A�����a�'���͈@�n�<9�Ě�h�D����Y�O��$hQv�<�ެ8^` pb�Umx��E�>�y�-��.`&��m��_��跁��y�jQ�j�4-84@�#~���-��yC�d]��.��4q͌��y���\��E�U;<s��0+԰�yBn���y��J23Yj��SJL��y��%bmP9�"H�#dX������yr�J�G�Ux�@G�D��b��0�y�h�9mv 	e��7jT��a˝��y��������'�/ǂq�q�
�y
� �\y���U:�%*R�G�!Z��"O���膽t7�� ��R�Y���A"O,���/ۇw��a�U�5A�p�i�"O ��A��} ��5i��q�"OH��a!W�^:�q6�8Z<Ո�"O�Y���X�pj
��	Z�i�"O�$�`P�[�QAA[�Q|a%"O�|�d���Zi��&�8��H(�"O\x*�O�o<bt���zT�2"OL� �����st-��N�>q3�"O��a3&8E�Fp��Φ8��1E"O����TP�����`k�<��dͿA��P�� �L�Z�ff[n�<!@%(/�v\�FȔ�E����oWF�<q7�R/��l����p=��i�A�<��_u
�I�� �mE��شɓH�<I���V ��d�4ZԶd��F�<�d*�%!5�r#P�a�&�E�<QƋ��՛doλ"T�@�{�<�S!��$1Џ4	[�=y��w�<ɷb�� ����B2]���H� t�<aQ�=��	$+�HP�H���l�<Y��� f <)* IO0P�ЉMg�<�T#܉J�씹'��Zl����f�<Qg�[���mqRB�~��)��g�<I!�?Aun�B���!g\��0�b�<)G
�#t\T������#"�G�<�RlG�V#�L�B��$�hx�2*�x�<1�6�*��ǝ "�q�ba�N�<��o�3hu0�Ba�!'D�p��b�<1�gX�V���$I�؁�T`�<��`Xw�:����*-rqƔ_�<���یB���k���|\��WěV�<A��Fv�n�(��"i�i�ƙT�<�@j���Hp��=NL:�F͎T�<I���]�L9rE<n�b�G�<a�b;�.���F5?�Xj6��C�<��Ґ'm��A�ƈ@]f�qV�K~�<�ѡ��R&�F9Z�t���c�<q3��D�j 
"큰b��L1�d�^�<a��V�K*����.r
��P��s�<���2J��I����f?��$�
r�<��i�uJͪej�)g�h�%S�<цǐ�&֌BG��.[���MM�<���;J�}R7l].h��=��JF�<Y�J �[Rxa �/�++���Q���F�<�@K�#9����ک|-RQ����g�<!Ӆڏg�R`��?O����%�x�<�WB	"�.�C�b�|F��EOE@�<������X0eo�(����P�<�ӂ_�2�:��.J�>�$6�L����'�`uA�lL9�ĉ���X!�'��y(#�M!E"��ĖNO:d��'cԌ0�Nv�h�a�5K+XYK�'��4˂DV5�X �0͍2�<�
�'����W��q�:�31�C��l��
�'��yE��&̀Q� a�"I����'���cs#�2N���E���(D)�'1H+uEJ>gRi�b�9*N�I
�'C��Rw�$]f>{��?,@�	�'z(�q�˽��p)t�Y� �r�j�'dAդY5<z���Ot3�mx�';�����ӵ[�:�˅�oz���'����Ƀ�8gb�R��vB�A�	��� MS��U"I0�x�5$H	|�"O��RU.�y�dC��μh{,����1lOe ��ϙJ���@�լ(oz� �"O��^S��h1]�o:�3�"O2�h���'N��Ц��M�詥"O����#�^��9c$�ͣ`Q��Rw"O�!�E[РȐ�)�]֚i��"O~�h���?,�"p7��S�\�3�"O�8��E
"T��1���c��Y�"O�I �^��.E� f´f��qѶ"Ol1�j��F@�@a$�A�j�3�"O	���н!�p�� �r���"Q"OP�`�3	�����l�z��"O���eH[ ��U#d�C�r�����"Of�(��` #�U��t"�"O�����7R��JrR�L����	�'r�K�
I96���� mE}z�	�'�&|z ��1�$I"@É/ep�J�'��Md��?ն�#� Z\
����'�\qRu�M�EV�-�ԨCTCr}q�'�V�)1^�. �A���I�"��'Πm� �I }BS�@�jJ�%Y�'0:|y�hS��2X�"L�`eX�'yT� D(h#���AB�.'fj�	�'��a5!�6�Ʊ# ��>#�X<)	�'�2�(�	�ޤ *���$"�����'�(t�a�I 	F ���0�p�K�'He�W">z��V�?P��,�ʓK�bH����q�|�'"<r&�ȓ�����Us�2�Qw_32�B�ȓ}&`aKaB�/ʸ���M;�FY��m~Ś"$�����3Kܱ9x�Ȅ�Z�6E�I�M� ��%î8�^��ȓ�V�٥�����Hv��)��ՅȓB�,D��ƈ:��L�@�Ck;�ل�
�̩ ��#�Ȕ��C�Q��`�ȓa�0,[���30ep�߄H�x5��!ص�w��:|��0�WY�V��ȓ(ڈ��M[_����U�"r����M�	SV��N.�T����&<�d<�ȓ"RZH����IX���*� &���ҍ�ҁ�;`�ɒB�Z�d��In� ת�������F!��D�и��X bHr0^�>�;�!��ZvTчȓ^ب�W�� I2�+�+[�ȓC(
r+C�Y�e���A1�(�ȓX���FlϦxu�|��+�
f�Ƅ��d~,���#F_�4 �EQ�-�E��=X.���28���&�K�����d�p���	|���a��(y���ȓ&^&���J�8���"μ)���ȓ7�.p����#9���Â\��b��ȓz3�5#v��(`h=)q�<O�T��(�Q�A .:��Z�
�v��ȓx�Q��Gf� N�gY�\�ȓ<�$��dD�'���G�E�f:��ȓ,Q<� (B{�.Ȼ�d��_<���S�Д�`<�˂ʲT��`�ȓoE�)	foN��zx��)�
@3�ȅȓ$��-pį���8���`Ո*aĨ��!���놵[���SG� �ȓ57`DRC�y3�+wN�4T���79��:c�T�?/8Y��_�q����EӣYZp����3Eg����S�? b!����>_PDS��[�$>�8�"Ox��i�<�(�C�	-l �H��"Oy�%���Y�B��%�P�+�"O�Es�
�l���#��k9J��"O�1{�*�R�9�D	ƫMAD!�$"O�KU ���s:R�2�"O$%c�O�U:Ę�C�
2�9 �"O<���e٥K0��LϟJ�H934"O��i1�A�1X���͌���r"O4�(�)�=8��+�6C=2�!��[Z�@}��u� �a D��!�N�+&�L:��Q�_�D� T�@�+�!��,
���$MM�.O��Y��d�!��%R�
�Af�+WI(����]g!�䗲��e�\+dh��[�!�I�^�N	���CW�X�r����!�$�I����V�|I;g '[�!��M��x-Y&�J����S�!�DT6/-<`P%�+B���*n��!�$�Ҝ��E&�<?s�X��MI>i�!��K� �:�h5��R<8�j��Q"o�!򄘥	��}yF
�=2�ށ� `��R�!�$Rڀ�F̂:|���p�O�{b!�dZ:~��gjͿq���Ro�#U!�dԒ*u(U8��S�u���S�D���!�X"z�����<�B��L��!�d��#(���%�Ô'�0]ʕ�]�!�:��`�ƥ67�2�q��T?�!��O9Wt��ל$�pk�c�&p!�D԰"�t�sl�w?�K���\�!��u��c��_�6)��d[�!�!��}�P(��V�ܲ��V&H�!� '�:i:���C��MЄi�4
�!�DV�+\ʘ��Ԏ*����')�56�!�ą(L�I�c��B�fuQWb�H�!�֙)}�%*�=v|�Ai� 
Q~!�d��j6�<��]�x�B�Ů�4!��_5C[6M(t��u���Q��|�!�D��~g��� ��d�(�:Q䅨S�!�d�C��<�7��kײ��5	�%dq!�Y�>A>��=U�B�r�ů*T!�1'G�qJkE�n��1f�tC!���%@�s����	�˜a;!���<M�r��4�׹d�� `��	�!�$��Wj��IX����ckT�6&!�I5���@Q�� a<��b!}�!�A��pR��G9ܨ9��o�!��A����S!�82=h)e!�$F�F��XJ4�Ef�|�����!��/���C-�ce�<�V�D�Q�!�O4BJ"�T%d��u��O�/!���4%� �n�^����ЬM,!�dM(��Q1j�u��-����{!�D��`�K&l��&��u�96�!�ę+oȐ��Aj�/�~MA6��*T`!���%�h��toy���s���K%!���2�B2�ߛ LD�I�(`!��O)	�v8څ�C�uEL�+7��y�!򤋥�q�*]�r. �"��(�!�J~�e�cƈG#֬�c�A>�!��jzY8�MO�O|�3���>�!�$΃/�������#�hQHG%O:;I!�Q4|6\)5k�-A~Le��cV�(Y!�$��u�6�0�T�RKI��CT<X4!�� ����m�)/�&��EP o���"O\��7-U2bb�!喞p	�"O�	����*5���ţI�ը�"O�� q�߸1������M�8zd��"Odq��$ǦL\Pd���K���"O	�a���k`QjSA�=�X�`�"O\-1�.�-h?��2 O#��@��"OT�7L�KF.H��n�<RT�"O���P�B8EC��ңN�Ya�T��"O~\�	O<�!����.Ig<�h�"Oxx��P����lӿEl���"O�Px0����`	�L)R�<S�"O�1�I��B���嚣��@Q�"O��u�B�#GLr�Ė6R�@�P"O�
WB +>���P"#�"=��*�"O�5[ m��4
w��>n4�b%"O���A�t�h���ֶw�{G"OH�SEɌ�H&�ݺ2
��x�"O��#p䁉fܠ�����W��p�Q"O"88��04�N�:��.#z����"Oru���R�"�`�Z!��[����t"O�)qŧ��>�I�@'Kǀ�I&"O��A�]�(ZF����m�N��7"OQqT�G��Q��	��ڄ��"O|:ecK�SYN�٤��m�24�7"O�<I�`W@n���JZ1�F�ab"O����L,xN~\���S9b!*�J�"Ol��4��������?~�M��"OX���;�$-�7	]U<��1"O�	꒣�.>�����>;�ִ
"O��s�)°��B�$�֌D"O^�b��V�A�z]�T��
s�h�"O��������U	7<��@'"O��Sȁ�4�>u��DUH�j�"OԐ����aRZe�ր�0��塠"On�
�����9j���b�|�Z "Oh����J3�m�%b
p�4"O�j��M��lY����:R���CW"O�<�ë�2���� -Xth��"Oĥ@��K���@F% ���"O\i�$�B�	��A	�n��@X�$�"O�@z��Z�.��%3���,�VA��"O 0+�FΦ6��y�XI��C��W�!�D�=�d�tե%�RX��oI�c,!��C;w0�!�nT�[Ɉ) �DQ>&!���r�h����
�bE�����k!򄚋Z8m�w��-`�^�yG�U�L!��@\��8��F'v�
i�'��!�$��j�¸k�gފJr���%�)>3!�$�������V�?dB�:�e(�!�$��°��s��l��Y��cX�!�D@��H�j�Aߌ���a�4)�!�d�$+ �ԎM.TيM+4���!��ϲA��pOZ�Y���)A)!�c�D�&BZK�����3q	!�$�d��f'�;@R|��!,�+!��E�Q���P�
�o�M�v�_�U!�߿r��p2�?�в���Hc!�D�	h�����W�G�U�R ޴c!��F�6�6��@�@�?��!��ć�BW!�/P���Pc���� � J��$��) d�3
� ^���#��J��y��̓Y�u����Yl� �����yr�]�a�&\�ƌų�`���޺�y
� �r�$NFV*��P75����Q"O����f/��蠤 �#n�
`�W"O>���MH'��ـ �9d^MÁ"O�i�b2S%<�/W�]n�l��"O\� �C�.Ą58B�f$)�"O"}S�kC0��n@m�`ezV"O��`�kR�]\���,ER�2@��"O*E�'OƉg��Jq���+���Qp"O�� uNB�T��
+
ּݻ�"O"�xT���{/D�XdKN�vB���"O� #��^�X!voF �K�"Oj���M�P�qc@�&�����"O���S�ׯ^���0�@D*6��Y�T"O�|�QCǇ$f���Bƀ>.��\�#"O8#7ϟ�Mؤ@��=Yx�D��"O�A�`���Q�`���)���h�"�"OD����K=]��E�H޳$�i�v"O"�zS!��n�Y�`ۮyd���T"O�#FJڦ	wҐq�NJh5�"O�EwaJ
'����È�nT���F"O��% ��$��c[�$D���U"O�d9�H�� 
6<�Â;c&�pk�"O�U �/�6��i[���{�dC`"O:y��FC0I���0��~���%"O����W7O?tPۡOW$�r�"OT%�EC6R��r$`x#"O@�;�L�06���]	!��U(D"O^d铫�--�tycŊ�8�l��"OX��*_�^J���M�X���K��yB�� nJ19'i�:8=�T�G��y� 8t`T��J��0�Ɛ�2O�8�yb�ƨ'ה"���"i�����!�y��*}���C�D�B�[qퟫ�y",H�U��v{��i�g�45tB�	K���D#�:�`Ը5�Z�RB䉞OY�쩱�U1����iC�+L�B�	�cp=b3�r�dy��wb�B��3g��Q��l��[#�B� _��H��(�~P���O�.�^C䉮I�8��jE����b��X/w��B�9:��ȧ`H$�X�����kOtB�&8y�Ѯ���x��Z��B䉔/%�����F�bqЦ��4�C�	�mQ��Z� ��*LL�� ��?�C�/[pu3Q)T#/�� ���!��A83��K���W� �����R:!��W� �����.4�^��Җ !�ߢd-ᒖ�M�Q� �8�b? !�D�9F�\͹!I��Q�P���G
%!���9�j#d�M~�1��R	BL!��Ú%J֑cV$�Iv����
РVK!��C7A�*i�rH9|qBУ2i��!%!��ϫ:�����j�/(`�3B�W2/�!�ĄdpJ���_�/ND	�4n�.�!�K�?��i{�[�5�~ Vl-�!��\�n�X<�G�}��p����Z!�$ٱH���a	�=�}1��
3 O!�dS�$�HԈ���PS�,J+_�~8!��.���� �P�bɎ�T!�䛜C٨Mp�^ ˔��'��7!!�d��r�x̈́�K�d0u�˪H!�Ě�ePy�b�ߕ���;��ԟ_�ў�ᓕX���X�-N/�D�7��/�B�ɳJ ��C�i�+]4%��L�u�C�)� ����]�V&��ƪN�]Uz!�"O`A�A(ŲC8b�b��-m^���"O��S�
�<7�p�h�%!V�]C�"O��aB%�@������<���	�"O>(��@�Zh} ��[�<�z�s�"O�)�D�R�$s$� ��֔zX@�0"O���b�e>��5B�Vxf���"O����9��g��.p|��V"Oj����O�a�H�%���s"O�)��'�p8�\�$���"O<pA��>}܋Ƣׯ2U��Bf"O�4*�F�&!�hA�aZ%w�2!�c"O�i�]//�t�3���/.n��"O����a�)0��`�Í3:�����"O�91ůqJ��T@ɭ.�d�8�"Oވ�6�%�jA�𠔢h�rX�u"O�*���i�&�;#O�KҀ�"O�BK!������bA�"O�m8K
!�ԍW�r�
���"O�󨞧Ov�0�M�-3�f(�"O~d�@A�%l��[Y�Z�Z�
��y®	�"���^Zp��@M��yB�\�i���rF �G�vY����y��*\w�̺a�Н-b�5�d∾�y�G	:N�ajs��������;/��B��2U��9Ҍ��8�L|�@�N��(B�	�<H�I���"�����7�B�	9o;������,a�)Ȳ ۟�B�+1���x2�Ä7�|}�(�b��B�ɝLx�!S h�zY�[�v4�B�I�#Y�q���9EҖ��QO�5��B�	XF���"�+y�Ω3��:Q�tB�	�-Bz��j�:4h�rmE�$;zC�ɈIk� 9�K��=�����Y�C�."O]��^2rD��s1��%$rvC�	�e�[�Ȟ<4S@�vĊ�/�B�	-N���V��Z�6i�"�N j�B�ɑ��i3*4.,�����*�PC�	�N�hm��'�}�����M��3BLC�5	�&@p7�H~���B�d<C�	�q���8�K� �hA�d�كh*��0?���A/8�*Ǩ&y��<@���x�<��jߞ ��q�.ϞI>�}yB��_�<��g�H� BpeY~��ò�JZ�<��J�<��
V���$���X�<����V��"���X�ڱ��y�<�Gɫa�Zh�uK�.ot��5)o�<1�C:G�$�g�֥��8��a�b�<��,�>h�Z9B��6zylL[��`�<i����;��E��8����"Z`�<��`˓4�N,R͞?c�l=2@J\�<9gH'N��� FZ;��!���FV�<	6턭g�.Mӄ�Ӹ���wn�P�<q�`��Q�����ebx�%�v�<A��R���IF�	&b^B��Ζr�<���A��4��I�c�J�`��S�<���D
4������!$ı(�-N�<�OB��g(��ak�@�XH�<�T�O`,�0��̓/�*8�e�B�<�"�
,����#ሖ�S+�}�<iC��'�|哇#��x!�h�y�<��̇�cn��#wJ�l0L�I��XP�<)E 2w*��t��h�a]J�<Y��R�?3��s�B�wƪ�@�I�<� �u�I�p��1Peƌ3�̱�"O.��' ����bD���j̓�"O�]0AK	��7�մ-^��ƛ|��)�5SD�Ѣ���Y��F9c�B��4HB��#'�sI��g��sbbB䉟m-؀�a�
��Z] �^|C�ɳ4�	2Cn�0Y�h����O�<$B�-[�Tt+�)R+WZ,�C��f�C�I(T�`�!'�6#�Eg@� VB�ɧ@h��06��r��8���BB�	�M�p`jr���0f�Um�p2�?i����tE�C��^$~��S��(&!�䎋M��l	Tn�,���A$!���U�A�KR5VKd�QS&��u!�I�3T ��i�.Y:V]	�GN���'�ў�>Ś ��76TI��!4���RGk+D�T��g�7#p����Y6_
�� �f(��,�SܧvJ�E«P�F��gɁ�
�*E�ȓe�Ub�CãS��:Ǝ�}-�,�ȓ#�6\0��D5j� 2B%�m)�-��G���7�J�:I��A#��^�(�ȓ4�i�O�9ʹ�Z��?�i���Lu�3�ս�`����{6��ȓr� ` ��B�a<�u�@���Mh��ȓ\�b!P�"3Xm�YH8Y� �ȓ"ެ t��5jc~��O�[|n��o@�I�w�Q']t�Y��,ԉ5�N�ȓde��2�+��*vhj�
�*k\��ȓ[@�daRF�/y���	NC?h&,�ȓV��!�َh�I��$�D���ȓ#���uFF2�������6�`��ȓD���Fl
6QR�eq��R�v���-c���Ď�o9���v@X����4�,�;T�� Wh�9ë�V$9�����R�ev�0Qq���-P4��ȓn]D9t�P2L&My��H�I�4��o�
�K����A�2B� +4܆ȓd|v0{뒻TP�0��!_���ȓu�<����Fh��o@@�b��ȓ38~����'g�L��М0�i��nj|�35^6=����&�!z�A�ȓF�v)�#� 
�Pl3҅��)$5��5�A��.Œ #v�Xa˿I���ȓ��+���2Rs��p#�<J���ȓe�1��O"3��q@�%�4ІȓZ{��u˃C��� !�	9)�\Յ�85zDT�P�60�!G��q�d���5K�HI���hZ�#cƲ��Єȓ1?ꔫ=���#�d�,E��ȓ&A�D�чKj$�M�*p����;�<jB�%���w���c*=�ȓI$8M��#�=4�|�!Үް��\��t�\�Gד<_�=qe�E/E�h��xM�Ҳ�r@H��G"=��܅ȓ,��@5�N�a�,��%Mm���f38��/�'�N� Ζ�Q���0�4��0�r�cs �	��$�(�	Qy��Ӭm�"�a7�ݴV�Q����:ua C䉄
%��1B	�Fu��H��Z�h3�B䉟}ђ|Ҁ�?[d��V�fԶB�I�%C�!��� �T�+ֱG�B�	�@���R�甊X8�0C@�{��B�n~��N��\�ʱ7C�=ێB�	#1�V�1c Þ#F���5�H���O����O�˓��� ��֥����W-�s��܀�"O��J�;e���#�*O��i��V����I�U0��ۍ?8q��[�7��C�	f�|a���)S�p��S�����C�Ɇ�E�m�� 6lJ ��\x�C�I m۸<9`hZ�w�+�
G��C��;0�"U�Y�R_��;��O�מ˓�?�O>�����01J"y��#�f�6���&ƞc�!��L�����)����D�[�y�!��#4B"�00x��֊�� !�$W�^���� �Z� �*<8�!�d�u]��b�cۂHnRE�P�M!!�䊰2�t9�	F`��K`H��!�d�TP�}A�n�+3^岵EQ
��Ip����f,:ҋ�hc�h�Eo�Xԩ�"O2�0aƙ	*щOB �Az�"OF�+p��y��<	En����P"O�1���0k�dI���ݼ(�L���"O �ҁ�����>u{5�d"O��28Ll�R��V`b�2�"On����@i��=��¢XN�@p�|��'�N5���mX%+�-�*W��;��x��ƬO�h�z���n�9SN��y���$
|\je��hK����F���y���74��PY�(�[{�łdȽ�y�IJ��1CG�� �f��t��1�y"4�4q#@IV�iP�[S���yB]�p�n$(�mK�a�U�<�hO��I�T�PRQ��.Űa����2>!���5/�	�aG�L�U[��.F!�d���6����rĲ�®��TM!�d�8*�U(s�-�x��3��70!�d]1U,�骃j(veBxӢC�5k!�䊲! ��M>U�䠀L�,^!�$Â>\6�ȠeK��xC�+�er!�D�10ze;��Xp�ڳ
�_!�dE�8^DkP�B5)¤���`��!�զ^1�pR�	�3�xqSM�'�!�DP)u��x���F�\ЩM\�A�!�ē�4���+y%p�Ap�)�!�$U�"���`mόtHy���2�!��znU��hΨY l��"X�ў��S[��0��,��=��Y
[�C�	�A�����0s��yǮƌx�6B�ɵ\� )o�60"�iJ�	Z	O"*B�5U�FP�4�P!!�\5y�l�J`C�I�H�b�����)mZ�$s �Ԡ\xC��.����g	
[�d��Cǋ�B�I�LdN�㣔<=�`�@j�	~��⟨�	B>�zfH6+l a�Jʧ��+�K+D��c��+v���h�?L���;��)D�A���3q���qb��a�3+=D�T���G����X3�C�$/>T���;D��؀@�f�2)��%�u��M0�9D�ءGa�ls�͊��M�_��$2D�\��͌P
|T�!nM2i"����"$D��"��KR��ZT��<f�� Kt�>D�����
fW&ئ��:9[B�Y �:D��9���ha0lQƧ�o>�0��4D���a%��7�����Y�����3D�Ly�jU@P�jE��ԃ�3D�Df�ΞF�d��gE��/�L i4D�th7�X7Kn���Q�Su�Hz�5D�X�0�C/��9���M|t��+1J=D�� �z��O�0�:	(2FD�8�4��"O(9���-4�I�kA�ً�]���	�wP��2a-��H$@��D4.��B�5��J@n�sG(9�1h&l'�B�	� �� ��!5�%�*��"����>?�C�k'֕��� >K�n��e�f���ΓN^P���_��-�'nYnѮ��OL��f�"��t�C���ȓZܕ�M#"І]��Y�~��'�^����#5�,Dq�$6���z#f�=�B��,(9�����m{�0 �<�B�Ɏ1��Xb� �	&��Q���B�	V�|�1#��/0$A"'Z�M�����J�Ik����/?Ē��W��4tZ#�[�{P��OȢ=�}��ńEM��9�7OZP�p�Ks�<��c��8Hb+>>���b�T�Y���OFV�:s�����h���|��P�'#�K0��-�V�� ��
�'���DJ\]^�q�c�?D���+
���?�f�4�l�)�ȼ3<��q�G����%�O�A�e��b�{����zjژ�P"OxL	  �"_z]����Ccj�"O�M�RÀqd����-Z���b��4���<çNk�h�ƤL�E�T���e(�5�ȓOt���� 1#G�Y17ON�C�Є�	��,�&��B `��7�Nf]�d��	ߟ�A��L?;%�4A!
8qPAu�|����Ei�
�*c��y�h��,0��h�'Z~��ĊG�
���"�pO�L8M>��r�;�M:2�ـ�.��/����	6��"<I`GJ6P�D��B֒ij�D]u�<	e��q��a3�ΐE'�(p#�Z�<�Š���<�cal�GP�%gi��<!�b	�V]^Xw�� 4��#�u�<م)F2k��+�O�c�,˵/qx� �';\AR���2|�,)�1C�>U|̙��hO?�)�"ٷ1(�1�gۈ1��1RG,^x�|Gx"��\j�Tq덣p���"�y��³jV����Dw������y�L Y3�����Fr % ��D	��x�̵P�*mC�M���&�R:3P�{r���W�]�*�E9!$�4SO!�ԛMYb���M���Rr� C)!�Ĉ�,�� �]9�e�G�$��9�?���~#)��_�IJg�	n�ARp�JU�<��ýD~0I��Y=��$���RX�<��h8OԸ���ָl��f.GWh<���Ɠ�tU���?o\�i�J��y�囜D���;�싞d�"eV�
��y���^�캄;U�*�25/��'�az"�!\���0�m��P��	��-ǽ�yIi��h�w� 5Kn03����yrK��vs�\1��ԎF�H��4�yb'ρ�%C�=R^T�A�gםe�T��I�<YD@�\�1(@��2$ap��r�[�<�w� �S��h�H��Q�(j]_�!���G|�X3g��P�����	A�!�S�cEԍ�� \�:��X�8*K1O�T���'a�����kTJ9Cd�.�����	��y�M��)Yj�B�����"�L�y��Bx��wDVE�Z��Ѩ˔�y��@���]C����괩�e �y2�^m�<
�c��#x�����?y�'�(5�ˏ�E�ؕ#e_�1o���� ���a� �FLBpC��}Dxt�����O,��I]w}n�G�Y�G���7�6)�!�$�
��k�k&[�xq	�� t!�$E(#��ܛRl��`����(ī)G!��؀"���"=n�y���3zU!�d��h~�m"���V^6u� %��\I!��@l�{��
K�bX+�ٌ(#��'���'�"S>��{̓8�,�A'L-Zw���U�N4aE�X�<�oQm~bl��K�0��D���CH�i�����]�T���y��)w�E�cƉ{Z�A��$�"�y��=����)��v�4Y#���y�&!R�D���D�N��-ƺ�y� �0�����Б����y���3>}&܂�8t�t��Rf$�?)���?)���?A*�J��?扰��a���6T��C�b���W�p������'��C�4�~	� �f�rʦ�9��˦�yr�Gq��P4�Ϸm&�@����yr�B�r�3�Jp������yR�,y��<w�nА(�%%؋�y�f��4�� �'�`�^"�
���y�+ K➍	�C�[���"DM���?���?I��?�-���d5�I�I�������o����0@�O�A*��O ����<n�
�g�b~�a�F�E�!�.~萬���ن1�r<`l�<X!�	q��(��aҽj�8���W!�Ě�"��q��.�� Xh�Cm]�uT�)�'M"f��ǌ=��iu�
 j���:
�'�����%Ej�asD�R�Ze�:
�'�� ���+T!~u{B�R(L`4j	�}��(ΓQ邰�7劻#U0��`g�%R��ȓk�mbԡG��, 4�	�6���1Q�,B�(�����oK�h�
��U̓#`�`a4(Eo.���Z��'cў�|�V�ĹX��� �x9���Wh�<9E.�	X��\@U劸;L ����`�<A���-W�h+v���<����#(KV���hO��;M�>P��N, �[���(���$����I2y��-�7
̫�v�pwm,n��B�I�|�\��!
�7T5��K�{��B�.!d"�r�����L�}]z�AVW�8�I~�S�O<�9�Ա����;#��s�'��kR%U�P��0i�0�D1�H>�	�H�fuR�φ�9�\����w��4��U���m���V�P��2 ԇȓg�Ƀ���|0f�Ce��,4�Q�ȓ<66%{�l�i�$I,Y�@�Ӈ6D��p����΄�(��ĕ���a�J�O2��&�)�'6�2I�k�8L�Huk�� (��3�'��h+q��o �5	`�D�o�Q��'a
���O��W��m�^ ��'2�Ia��O�I��,W.�:G�-�N>����)��OU��i7�1��h�!��ҎD�����+N�����#�0?�*OL�3DE-I}���F%ǋOI9JCL�O��D!�)�'IF��4h}�DDx4*�#VLs�'
���ꏍM�^�z�D	�A�ij�'�f�3�Wd�*�i�陰}@
�{�'��!���	u|�s�Ҁq���J>���IWtv�+@�N�vp����(!��@�In��Bk"`pؕ��C$!��f�(�z �H75�]�� C�}kўL��ɥO��p��d����#��(:�B�I!2�pq!Ge�(p�<x{Q���o��B�	4")�g)<�(�1E�kvB�)� 
ڡ�|���JC��9���қ|��)�9�v�9�,]�q���I�#�C�	\���#$b�1��t��ә��B�	���A2��R�o�n4[�	<C�B��.\x@�Q@�*t��b�-~��C��'2����h��z}J�K�.�JavC��5	.�Q'�E�\�(��@��	FVJC��2qs�(8��~{DUC��+lbC����ᯃ�)���!�&�!w# C�	�wCbѢWӌ\��4�v��#RUB��sB$ t�?v�ii�FӛFq�B�+۴��g��qЌY�O�B�#E�h4 �B���L�fgLi�C�d�Yw�в(�6��Fc�=%��C䉣A`\���"LtD��@$^#)E�C�	�{Y�l��O�(	.����F��C䉿
J���l�0\t���!�!��C�	��f�� Oļ[7@5��AȰG�jB䉜B����Y18 q0����/J
B�I�`�y�4ŉ:9! ��!��q��C䉥n�E��%��b���ɀ�tC�I� D8��-1ڵ�A�44��B��%p���^�zn�C򋛨v�jB�I)>BL�qf�A'TE��@��>k�B��9\{|A�� �#
]�1 ���f�dB䉀U��y�GnվD����R�@�B�I�Q����MP� �Q2�E$#���'�2�'n���G�eE�q�%-U�IK\�!
�'�Q[�cE >K��C��6VOB���'�q��a' ftaB��ѻ7N�(C�'4yX�D�6�訂��:Ԍ��'�����0g=���ǜ>9�|1 	�'����o=�Q�B��,mtT��2�'=ax	E�R��yuK)�z4�cOȑ���O0��ă������A5c{��j�$^	�!�@>���)�!tT���-m�!������C�%oGy�ը��N�!��,xT��;G講��ˠH�!��<A)�q'� 1

�
rĘ��!�1z\P���u�Τ��)"�'^��c�,)7�C�Kx9��ە2*�p��"D��H+�F��ic_�;[D�r��=D�����QG��1�"��q���'D��S ��=	���h6G%an����K&D�(X#"H�\hK��{�8х+(D�,y����F�|�"F'�F2@�0GC+D��9aMܘf��!�uL�+
.�jg=���Op���L>~_f�3�'�zd�U�WQ�!�iM�� ��ژ�@��"y!��(!�Vy�CLF�B�L�k�F�oY!�Sr�`��@�2��%�@��Gj!�1�k�$�ڄ[e�Q!�D^87
�$#��_.X��K�dG�\!�$͸0&��#� �꼁JU�ƻ`!�Đ1A-��*R-�ح��"Ąy�!�]F���䊞=O�V�[k¬�ȓLh)��A�G���1�%���0�s�L�	��@9�B�1<ц�LԹZc��,d�Ykק�0r�Rl�ȓ]�(��+�=��HK��̑��D7Z۴�Y�qT��� B�,r ���i�n�Ӷ�E� �Љ#�^?%Kt���(�|��&��� ���r�ʷ�}�ȓ(1,�`�Gݑ8v��B��YA���S�? �����9�#�J(FrƝJ�"O�K2��2�x�j@�[�����"Ob\�n�{��<[uH ��L=(c�|��)�Әo��Hے�'v�� �7�ܼMB�C��2%�z�2�d�7 !�B�k��
%NC�	�$(B]���J�i,�zQ�k�C��;S���qE�U�1K�b�u�C�)�T`cU���0���V�~�(B�I�vc��@�J�?@�6y�ÊTSG^C�	.�~�↓"H����d��!u/C�I=1,ua���9��x�ʊ�>c�B�	�H��dо���Y���%�B�	�WaB��C�84��x��oƧYmbB䉾&{�c�Z+� �����dC䉿0Wh�3I�
fʪPb	�,(mC�	�a���M،an�D�e�F�e��B�ɑ6��a1W��?,a�H�$䄺\��B�I�H�X��>m�&�ZЬA1�bB�	?G�ȉr%^9}�L%�Iˠd�*��?����
<݊yP�	�6��-Z���!�d6Z�r����:�:Ã#8s!�D@a'�s��L��!a�׊g�!�䆯h�D�[�
ǅH��q[F�9N!��ɘ�"�����j�3���9�!��ή���(�*]�q���+�P8 �!�ā8n��y�BW�IJt������_��Ify��i8f��݂�`L�F(�5��wk"B�I��섘 �ǩ�<|)�_>;ܴB�	mR�����GB/0�:�/�:Y�C�I�^F��v H����J�hx�C�	�-�D8�g�R����I�J�\B�ɝu��ݺ���G[(��甆0�0B�	4P�4�u�ɥHQX'�������O��I�zL�̹��=H�����kR7R��B�ɋ_�ڤb�	�eD�Q��h,�B�	!u���j��V&	����N�[;6B䉫#��pIA���%NP��Ƀ|'nB�&hD x���<2��Z�i	�U��B䉢Cv��0����C@#i,�B��.,1j�)���yY.�i�� �O�X�=i���'�d޹W`:@)��	&]{tpȒ�:u!bO�2��w�E��.���V"O���ƃ��!��e�4���T1"O\e�'�$Y��Tf��@�R �v"O���K�+s��������}h�"O�Z$fA.$�U�.x���"O���s" e�֙z��w �W�'��D�$ضI�hM	{����1��	i��$���2�h�yV�[a�xc�':D���ƪu�����{�8�q@c;D�lᑌ�`��S�lY �{R=D���@k;N�� ���54⮕8��:D�T����  FX�d�E�!̮���&D��x1�S/��۶ ��Q]���F!'D�\@����RP�c����ur@�#D�L�Tk�r���GM� 5=�87j?D�t���:U� �L�7��R��8D�ԙ`�#-�|P�R�Z��P��8D�hr� Y#~*��e�#G�t��4D�d3��R8)�xM��C�PL|@ɰ�3D��KU/�=/b�����"�J\s��3D��1�陛[�h��4$�Q8���1D��ȑ%��}O�bD�'J;.h��	0D��`���,t�s�6DX��*D�� ��̘�GT�Y&`Ob���"O(�cr �qPd!Hf���F���"O�$�D����.��-Ҁ�� �"O*�"�ǳF���H��9]z��7�|r�'ݶ�&כut�!��
3/��}[�'�j����e��� � 5A���'��0�Ď(
3�|�plI�_lD���'F�3��a�����Ԫ�0�',H"���%  T�`tM����U{�'y��#7k6���*g�јF���'9ؔ�5�٦_������7@q������?�����O�b����ߕm�v��2
2-��32&�O C�ɛv�B�k�'� 1 l36mM�rC�	�|�0��gN >��Ԫ��_|�
B���ha!'ɀ?G�ΰ�'��{��C�I�lsz���=a`�B�g� }DB�ɕp�4�j��E�0��_=tC�I+��|�!�?�lܣB���!:��$�O0�=y����6�2����t�3�`��y�xR.O���#�O�i�`�� �4ѱ���`�x��0"Oh�j�MӗM��Q���3�d͡"O6=�Ѩ�8+N �y�F� 0Ѭ��'"O�d���9��Љ��V�PI�"O
dS�+B����e��&s�r 	��'W�	7s��@��`p�W	�L�C�	6Gnx@���N��@Jչ{�&�O����M�dǨ����F	��Dҧ���ll!��_�T��Řwˊ1;�5	��	�%i!��`0��B@f� P�4�r����$U!�Y]�!���j4@�e�F�!�$K�VL~Y�eAϞe�0�H����{��'k��
s�������/�����SX"C�ə#ǲhpw&U�:���D���C�4�B|j#�Z��1�"�Y4�C䉅:S�əvݕG�z� �"ׂ��C�I.W�rx��D*%Ԩ�2B*�/Z�LB�I�L�j��F�Y�](�L��,�tB�I�q���㑄N�%����Ҟ4ŀ��$�O���1�ʡ��F&���B&� B䉦%�L�x�_=q,��Z K�&y��B�+*��$���@+T}iA�^	WnB��yh�pJ�	gUJ�;a[�.�B�I�h�҄B@�JVF�x2�W*{�nB�ɨ�*;ĩʈ����#U�`M0B�	2U[�uS�m�51�9PE� "m@��De�H:A쟕p�b}J4�޳:�l( i4�I[x�x:�͋6	�Lӌ;|�1R�~�<����C4��	#ϒ�yR@���+�}�<�ǎ�v���[�,ɑ��y�<���ҧrr�,a�l�q�Ҭ�t�<���C�	�R�A�AP�u�me�\�<���#"�d��5	]��EI@X�'a�d���Z`�P��P�A�\mH����x�$դe�`A8�ա`o�И�*��!��/Qf�õ�:�j�����PyR�n����@��<t%S2��y" ��ΐ�S�fd�¤
�yR��*�t--4����U�4J����'xN���.+d�< j%E����	��?i�'��m�!i���ٙ�10���"�rو�n �B(�P`T�}�r����'��	V�� �K�M:���ѣ./ٔ�:�A4D�$Vz3��2�BBJ�^)	�l�M�<���»:L�bW�AO���"-H�<� ��B�o�x�z���jԬQ"O ���a�J}� ��.T�ps&�':ў�_�'^Q�!�~ ɉe�
$�A��'�Q��FčU:����	R�*-O�����$x�0��԰a�fb��S�_t C�Ɏ^�2��Hn *0���F�S"�C䉴*�Q���$[eе���	�K��C�ɑEY�\XϚ����$$��lC�	5VCj�S���Րa6�A�����D)扢b3:�z�&R,_3N��#��4k�B��E0TV�ȔD��ec���"-�dB��.ض)^�:�I0�?Z�&B�ɋ2̪4�r�Ep��ӯ̫Yj�B�YX�@��G�$J1�)S�܀;ɆB�I/�H���;%U����Y)T�@C�	!1��@�P�TY�-�sBE�i X���OV�`�p��#��a��I�1 M�T�ԇȓ4�L56Gϣ}�ZU{�^-$�α���B<񖩓�<��2�#Q�1��e�ȓ8�䵙�-�^���@"��Hj�y��6�@02���!���j��سy�� �����5�ƶ8t2�O��Y���ȓ�	��M�+�.x��N�b�N̄ȓ���@&�S�r�i�&� ���5E(LHS�I_�<�ǶB�б���Ʃ#R�ߠI>�#�	n}����V�D��KД��T��g�ą�nd�,���/�x	���5|��ȓ)�nmW#��H��h���9N@��f+�E�p�:�H�8��˹a��هȓ ��q(R�d�t�BG��v9�h��h	�ѳ��F� 6(��D�q���$�h(�֙q��s���1W:@�����o�=~��d'"X1]$���hȎ�S�h���A�h0O��ȓTt�1�C�S��e�"H_�9�"�ȓj�R���1����%��9��x�ȓs�±�J�i�dY:C��;9$��R��@�E�Iy�>	�AF�d$�ȓ#=��AcQtᰍ�vKR�%���ȓ11@R�[�r�(�I����2�>͆ȓ�(a�Dv�I�'Ð� �ȓ$4R��@���+jl�Ӣ��Nߔt��apM�'�� [}����h�|I��D��)�֧�(C�J�I`���pe���O�ⅻw�Ii�h+��N8%�B��ȓ%ӊ��֩/8D�S���f�:��� �yI'D��4���u-�S�ԅȓ�H�)���Њ7.\�n��܇�)��%0�(�7?����#�\�Ll�ȓU�>����s<���Oʃ1a�m�ȓ,��Ah�ė��&* چ,t���'�~�;��ǫ4�Y��Đ��h�ȓr�0�Br�S�Li��	|���=[�[4�řp�(2��3�i�ȓ0��<QQ`�JՠrDj�z@�ȓ��hf�P��,��II2�9�ȓ/*��Ƣ�:=�4DA�oZ�
>d��x��d	� ܰ!v���&�Q$e{,��w�rI�Vj^�N@V�P�*H�+74���Bf$�-޼[��*vE�QJ���b�fM�4�13s��c�ƓF"�ȓh�6Q�G�� O4�4a�- ���f�
�p&�F
�ۀ��@�(P��S�? ���
� K��Q��Y�0� s�"O豲SL\���E�V1l�옪 "OIۇ	��$C� K3k�P�H5�"O&�EJ�&|CL�rt�ڳ+sfʣ"O
� ����F��FI�E���"OP����< ���H�3|h "O��{��	�R��s�ϠiWd<
"Ob�(�	
0��5P�i[�b?��A�"OV����<Q�,ڲa�|1ؔy"O�mԢ��0@�[�h�>��š2D�T��!��B��@��\!*8�g�1D�Zч!C�BI7������'�0D���5'F��!�g�NP�x%�/D�LѠ��h��K� �xh�B�0D�9AJ��>�j��c��V���r��:D�P���H��{���]=����-D�{@�*εy�GÕny�	�.)D� scF�s��a)���>d,h�u�%D���$�	 *E5�5F<���#$D��r� [0cO�{p�θtl���!$D�4����F�8�b���CV��Di>D���ŧG	r#Pd�,KO�\� �7D�\��DF!r�;&�Iw�R\(�7D�$3�=:(�h�/�/3�Jla"3D� (IW-z�|u����6QwJ��6D�P�䁌~��DF��P9�R�6D��;!H�%!����v��A�2yI��2D���S�4jvB�Ӎ�LOj���b%D�캆��$M`�/E�f9��K�i(D�<UJ�!�
QC�@�?~���'D�D�$/�4]�²��C������'D��1�ɹ�2t�b+_x�tH��1D��2"G�(y�H�.x@./D���A&�Z�Ӭ�,�p�jFJ-D��� '_8|�(��cH3X_�k��)D���q�}�!���!I��,
�4D�,)d)�'s�jU#夃�}:�0S3D��j�eu�P�W�.\^�I�5D�ly�-�jE�A�B ���3D��V�+	ۄ5�Db�Z{��AH-D��a�N�m�0�z�@�u$J��U�,D���#d.`f�@K�bʂ�*G�)D����IQ�P1ࠨ����(��a'D�X����)LɀD�V�I(�8D���&�6R%�},�Q�$D�<{��L�4]���D�I>�
|��d&D��`$��
7�䩑�Fɩ��y�p�>D�<���,���#/F�s]����.D���0oQj�s���#@ԥa2�*D���Ù�A9�j�|Hv����)D���V�� K~d�P��y��rp=D���$�-t ��b�>C��*a�-D�(�!��
	(}�� �T���!�$ D�$�H�cК�1t�	|�D}�1� D�䊃��Tk&u��K�*��9D�xY�g�4��h�Aj�@�)=D�Y��>���nC?:Ƹ�1�9D�Ȋ�L0 lr���b����g9D��8���n���rrl�&T:<�gH"D��a�	EV~�P6�ɪ^�"�r "D�P f�	S�D�Cb#F�I,��SE� D�x�!FõR�V=j��W�a����;D�ȹ�aȰU4���-�TO�!���9D�pjr��d���/X%4)�X��*D�� �{��T	�e�ե@�!��9#"O�UA�L$VT����}��"O���`-�1]�����ɸ�p@��"O2`�U�:m� bC�9պ���"O��HC�S������M�$�jj`"O0��u��=�T�	���11�:��"O  ���=�>�҂�M&2�ZD�d"O�%)�=���B��׵����"O4��Uh12f����W���Q"O�0��� L���`�E�9g =�"O����V�fXa`�V,8p�-��"Ot���A�)
���Ϟ�a}h6"O��	Q�7����M�*~J���"O�I���Ñ|�T\��坷HFR��F"Oh�nK,�80��d7�j�"O� c������$��;\�1�p"O���ve�<qjYkw.X2z�a"O$�I�6 ��P.$�=3"O�RA�o����G-�|�R�"OtLs�M>:��I�"�\���f"O��B�I�#T���g�Y �ҁW"OY�Ī�3�j�r����1�<i�"O�L1f?E$�� �C�"5K�3�y­H_��M�z�-Kq�G+�yBA-D��+��қs_���0���yR#��*��+o[��M�yrB�-\����l��gలg�=�yr� f���@�[nl�ɵ�ē�yo�u��͈p/˂iD����H�yRおoB  cȡw �<���y"��?YCZ\
W�oh�)B� ���y����*�Ta�G#A�m���6J��yr��{ݢU!��D�bx��Y��y��ѕ\F���϶=|���A!��yb�K�ހh��U�mج�y"��5\��c�X�-���c���"�y�.L0ʸٳPW����c�3�y�
wm	`L���p`-�>�yB�]�GL�𰐥�)E3a�N��y2�ۇfw޸��僥59>l;��I:�yb(L5B�l���^�z�*��GfϤ�y�+@3{V�R��!H�diR�[��y"MD0B���R�]�	~6���)�y"�ê�ڭJf���k�e3gO��y"���s��ͻa�J�y/��Jƀ�!�y��ӯ#�4�PI�8F�HUH�Þ��y�C����aA��D!9�R��t���y�� @����&�ս*༒�N��yb�Ǘ4��9� Y� )��(G���y���&����c�@���q�F�"D�0p3ELH#�
�f�)*��I{D,�>)���ӑ[�~�1��Q�[d���F�#��C���{u��@�bd+�-��ݬC�;XG��CcHE%c��
Sϖ�#��C�Ii�.t+2��4k���#��N^C�I�P��1�m�R��=��W���C�[�t�P,�^���4H�
-m�#=9��T?�Z5eO�q�q��)I�zz`+3�<D�����!5����O¹
蒥���f�~�=E��4b9��kǧc2�2@��b�8�ȓk�>��ni�ÌO�z����I�{��q%�4��%�'L�&�؄�@�qd�C䉫YGd	�B�:)8�K�q��<��+�ȟ` ��LǼU+�PYq/��d@�ܺv"O� t�q4�[	#A�I"!)D#2�0�BJ���|�?E���s
d�#�W�G��t@e�\��(���	o~�	�U�-�W��:\�lԁ�鞭�y�m����-��(qYF���(O`tç:$�A���-�t���ht���	|~�h��nU���b`�	8�fY��Ӕ��dLs��ywfE�]�$� �Z�DMV  1%G��hO����&&��M8�:#���0g�ܧ$'��b�����`J-ܑ!!��s�u��.�OO}�%����f�jč��l�؅���O(8���*[�\�3��$���@��C��1L@��҅N�y�C��_-$��C䉸<�aWi���pBݖ��C�ɩU�V�CbD�'9ܝ�Z�E*�C�I	x�a��oT�k]�H*P�$]��"O޽�2A]R&����_�5{,�1�"ObE�#δe�a!����&dB`��"O����@��Y��츁%J"�jMK��� �S�S� �b�ɞ�H1��_��C��3�Z9�w	�� �$�j!����<��l�p��ɘ"H��Ez2�_ {��9��fd�fFǫ�������Xl�ȓW���"��C��E˗�G<2����I~?�L>��ۻbq4�ᫍ�K�Y�SH�z�<����6I���	@�?Bs��Z׮�s�	��ē�?����Ӻ{�Λ;&��WE�A�P2��x�<�D�T"%T��J�	��cb�[�<	qJ �*܎9iB�������@W�<)t��8Q*�2��7�Q�2��B>�'��{  8��6M�!n��l�&��-r!�M�� ֢!z"���ɺ#��qBV�<iv�׎"�U��K��+��R�N�<����m��D7��u]�c�N�<Q��<U�~� 0,�V�*�I�u��p=��*n^��#�"�W�{�"4��Z�d�/��Ov�P F@Ep&�9�S�Ow����"U�Dv�L�ߐ����'Q����%C�.��d��D���T ���8O�@X��L367@�I�.A/C|B͛��'n�v�	"�$�'��Y�(�2z h#�"O.��`�$yJ�)t=��DX�t�	O�oQ>��qO�=E��9�1�<�@Ԫ�M<�	F����re5`��R�x0�����1#�ʓnIx�5��������;Yr5�ǎM2Y�Y�Dː.�a{2�D9Zj0y!	�5skD]���^�HM��&����	�x�(��5/^���C��Q}K���$��M��Ƈ}�X�ԇF7ON�,z��I�<Q#gP
gf��jC`�,(� r ̅D�x���� �?�49óN��N�0��c"�.�'ў�>!�V�Қq\�t����m�N0�8D����MSA�)8�APY��l9T'7�I�y�鉒("���f�F]��i�F.h���̟x�4/��)���h��ʧ~ޔ���!��nڤs��0�qhE�|���B�v��B�`B��	V#:'�\4CĈ�+'�^C�itp��]�m.��$.ܽ!�n(�ȓ6�1��4n�Y`�@�0Qr��ȓfW��)@�˝z� ��6�B�#�&݅ȓ{"���tVv�k��E��u�ȓF����B�S|���I�|����ȓ1x���Pǂ@Ը���'@M�L��M&(�nS�~���ej�/}�!G|B���,}X^�lX�#�a�I>C䉸	�Ճ4DN*}!u��.�
�B�)� ��ҧA�'����� (J��j1"ON\�QD��䠼T℔1
}	�"O��1��&@��*�Ι+g,&�Ca"Oh��M�=�`�C��!p1�"O��J1 �`��}�4�q�D�rV+'D�(��/!\LAzq*����/$��X���I�*:� ̑Af��n�����A���	T��h��B iN�=��]K�f�"6���}�D>�6:6^CG�Ž0��@ЀA�)n�C�I��4 ���,`���L�%d|�#<��j&)@EAݟO-��I7�B�lݠ7�'��O�Q8�&h0�)�7(ĉO���^���'#�曟�m�X��#n�UY2*
k��) #͑�	�D���r�j�C��C���ē�+�,�]d�I��\��}��)�)PѰ���J�ȑ�L_�",qO��=%?�"TbעT/N9����SE�m��h)�[���=�fʁ{>śq�)�V �#)�Z�<y�D[#�)p�	
�j�G~�<�b)V�dxp����ҍ��:��R�'�D~���>�;f��h�D&۠k�D���'(5���M�{�A��ΛD�F�(�JN�s=��$�<E{����@�:�x�A�س�Q�O�yr(R�h��Q��荐I�f8�b��y��
�@��mY:6����ƽ�y�l	�fY^�#��L39~�d�Jׄ�y���Gw�X{ Q���I�w%���<�����"8�&@.�$���m��9!�ژY�Faqa��u��<��.�:Z�'��d5�	f̓P�PC��QIl��/D:^̄ �?!K�HD�Ĭ��p5y���C��x!�O��y�㔹(S��
���m߄)�7ᅬ�hO����/��y�����2�Uz%�K;!�d��{��p�MZ�8�h���D�0!�$E':a�	a�+T�=�R��fOJ�r&a|�|/��(��!���Uw���AI�.���CX�� �/zj�p7�Q�c�x�p(<�hO��)O�ՠ5��C��p{�k�"*F�C�	:R����ƈ��-LAc�Շ/��C�	���R��0���9�!�3m��C��-\mB�Q���3m���#T7�C䉴R`(�3&ϩ �����:0�C�I
����$��~i��e�c����W	i7�5=$��fen�OP�=�}��
�}��D%�AU�&*�u�<�"`#t�౺���S,�[QaOt�<!!�Ns9�:�ݙe�}SfZp�<)���=S.� �����0�g�n�<1fݞY� �Q�j�rx�f�Cm؟���k����d }�h �%gg�O^��D).�BX*��	�|pq���^9?�a}H6?9�Gƙw��m�ᧈ>&��Ey�<�g(�>yY��S���o�t�<3ʁ�#"]/J~V��#�Dp�<��J�;��d�b'ܳb�\��h�<I�/D*^�8`�.�3�d�F��N�<Ʌ&��!ȱ���L�ĩе��L�<���+��ע��f��[w�UA�<�G)�P���Ə�k5��kwF@�<�3 R�j*�|[��;r���af	�B�<��/�*Ծ��� �5eD�x�THF�<I����($��I�/ӱi'Ld��@l�<Yv�܂u��d@$��i)�I"H�e�<I�Ӵ{H
��)�,Rm�@�E.V�<9Qoاu� �+�B]�e����&[�<� ʬsVI $��x�nB)�aap"O>b� F�^!W1|n
Ty�"O�IV��)���	�jˌ���Pc"O���1�B�L1^�Wi߉<~�u��"Op%���&N��Y�"X�'e&�9�"O�q�#�&�Y�a�9s���A"O�l�"�ͥv�.8�Eƅ �j|�4"O��u�Q�@��$�aj�Xz�"O�@1�K�LaΈ
v�� t@�M�"O	R�ĝ?�D���݋C�	�"Oِ.��~��-J�'�:UF
�"O:�z��ĮL���%�BD��"O�I�v��$g�22C&N_B��*"Oд겢��>�Hؒdj�2\,D���"O��Y�"�h��J�~!�"O`��ТV'�p(��HԖx���9�"On\�r���lE8���	loެ��"O� �fKȟ&�"hI�	�iP��"O@ؘW�� 1�`BU7)n�q�p"OB�B��ª#�F�����)��y b"Oh��F����x�� �!��`Y�"O����X7"�\�8E ��^1jA`r��q��$��d[����#ˇ�CP�I�8Ӝm@�		%���h@��Lh�B䉉vZ1�W�<���"� ��2,hC�ɨ��)IE,�kӐi���.3�"C�I�;�t͢��_	;�du��L�DC�	1K4���KZQ����
v�B��$(���@gD�7Z� �
C��C䉒z.�\��G�#GH��.ҽpZ�C�ɝC�*@R�D�4|�l|��>K�B�I"l�6�X5�,Wq�X�c�Զ��B��1��H����y���"U�,��B�	5���"uO�Eu2�0�,c�B䉯HKT�!NM�4�D�)�[�jB�	ks*q��D�y\�!X�u�zB�		O�����e�9*bœ���C�ɠ���� ��H�]p��S$z�C�I�G,T`�*.�I�*Í]�C�	�A��r�ƻ<��)�.��1�8B�	�*Kؼ[��B�"��:׈U�"�B�	=:�>lv�_�5��4i�4tI
C�5yf�2r�DS����A�){Z8C�=?\b���a���"�ϱ��C�9�<�Ao#F��J ��8�C�ɪRe��b���Ԩ0�-�0m!C�	��T@���]$��(E6R<�B�I$F��"�,�V3d<�S
C�k�B��$�t�	�IW!8J���gM����B�+r��l���3���j��/C��B�I�4�L!0���V�` �a�)�B�+���.�(��}����hːB䉡�^m��Ȗ)7Kp}�Ҁ׋�JB�IQ���Z��H'�Vmj��^@��B�i�VD�H�n��QƆ6,C�ɉ'I�A�',�p�P�Ʃj7�B�I
\e���LJ&�.�X�&Gg��B�	��΀�UaV�¬��_�@H�U@0D��@�ώ	\�ڈ��X�q�p��=D�pۤ�@�Q��B��զ�2"J�<�cτG�X�� C=z,R#UG�'@l��)G^�OL�u��
�c h�nF�Rې�[�'�h�C��&OL��g*��V�%�kV�3C��{J>���OL�׈@�9[���Θ�Q���z"O��X #��x@5̐�xZ\!��i	�3�d�
����)� �=���8=����Vl�#SPX}cQ�'҄%)�j�(j&�=�� �x��d�m��3u��B�I�I�z%`�O����q���6��b���DL� r8����S3o}B�abU�14���q�,ZB�(dv���\�A�^,�㫊,4�:�g�=e��O`D��O��b@΍�	~��P���@=��:"O�`
�F?I3��T	�2j<8�i"� ���e�$M��Ƀ.�
���HQ%n'd���۽z�t����-]Rvu�'o֯�?!�*��	*Ł����P���m+�y���{j���`��n��5�܊��'�@�CQl��?k�T�J����C�y>@�+7D�v杈DVXZPb��70�yf�#D�����܌:.�9�i�4MFe*6�5D��y��Ŗj���
�mB��F�C�<D�0R��ͨ-3F�zG(T8z�UqA�6D�$ TJ�,+Ȃ pd�I�Ne���6D�P ��)�P��&)MA*�s�3D�A7�4o����P�؛L0��SG$D��h�/��*� �_u�:BfP�㞘��<Qs&�(�(�'oE�1/l(�� 
7d�X���O��rO��e���bA��3k�kA�V.f��UA��˪��>	 n¼ �� �'�%" 8DCp�Ƥ �,�3+�`�'�� �$��$ $0H[P���<�0M|}d[����E�\�U�n���>;Ȍ9�Ov`��ʈ�1+�\�� ̘g� �	���� '3���C�Ǐ-XE�ċ -'(����_��M�sb���'���A�"�K>-a�Ɉ�:4vD�gL��/��5�B$�%����ԟ����(BLb>c���g6�@gԃj%�A� A�#�~�L���s�2��,�<x�f!��
��Ȁ��`��12�ջ'ln�~p�l���=aS�^!FW�����Bq��:d-O$67�	Z%AP�@��08�o�\�����Joj��!��h5M��i^������*u�����3;<v�')°h���/��yKo�4+�O�u�f@
�|2�X�fT KV��~���R2ψ�SLY)��)2G��D�_�2C�	M]��Sđ,Om�]�dO^':#�����Ћ<J鲴�޴K��a�S���*P����l�/3��Y��J-���G�?�\Y������џ�;�D����cu1OHdJF?}+�̂�Z�.�F�S�(O�W�ZU�"�/?|�y��T9'��<i��'��`P��҆Sږ+���`�Q.O~\9�(ڬu�jd��'R��ġF���z��5m�%c��X-�� U�J�MD����aY/T������O���$UaCF��3�.0�<93v[LX=�>���:�+�0`d�dT�bFJ��C.N/1�2-s��^K���~�����ؔg���9�ʛ�
!�2b؄{��KGq���P�Y,\v��4�8D}��qp�����ҵ�x����ݠ;�����h���V�_��A����u,�"vS�i�҉���O䃗jֲ"��Y1�'��hpN�=�^\[��LJ��yC��S1>5B]��D6#����d�5E&=�3�9�Fl;���X��|��@ޕ5������ۘW��-zQ��ӷˆ�la�DRud���޿^4�h+�*�n(8I�!�g�PAI��ߙ!��M�0��s��(�����>A�h��`�<0�ƪ�5X�`����~���6T�ȥ� �)K�@�B�L�a�|3�ȝت������$O#m$41�-"J�R�e��k<�פ�@��9����1�D�v���qt��,��h���'�R�8�Ν@��1�*���Q8=p�n�UV83�,�����R)8<�����x4�Oڥ� 0j�Tq�a״�tA�JQo@$��	U�>~AC���G��00�E1i�ZmGz��D�2=B��8#��b吘�p<��H�3(ꘘc뉔Bc�a����R} ��7K�g�� C'�čC��UG�z���`�[���#��V�Z9Ĥ!w��+��$��1W��
*���%-=<h�Ń��q���2Z?��q�	
>�M+boM�.�| ��m-D�(S��V�q<L�0�DIdXr�8&�Ȳu�l�.ʸ�B1�Ƒ����(�w��9��d�Y�>���@T`I�'��ՠс�#���@�]�8�h��o�:8&��p'��h�D|���d� ,  �.��\�D���ygF"n�$��-F�'�X]��CY��~��'Aް�1h.�L�Y2�a���CY�k�ry�}��x��Ol2�c ��%ɶL�E��-�Px҇�7!��9X%���]�|��ǂ*9��� ��C�y{r�Z�~��Ŝa��q���w�l���l@��p<!$������&?�m}K*��gD3H~��=�T�٧�"���,D��vd���R���0�x�@#}�E�� j"����O`.��π �8��ʒ�74��T�!=�y��O>�i�NY�x�f��_�l( �*� P�ɇm��I44��2`�3�s�26��ż+��X�4�r�b��QV
�3Wo(<AV睩 �T5 �e��k0���D�5m�n�2-��M{`-&?����L>�'T6�;r��	fE��D뒛M!̠�	�ς2�OΤ�'��]��i�}��蘔j�6D"���hO?娀I�:&� D�Ī��'�� ru�e�%�E�i�AQ$�f���
�`6gs��  �<�
�E�R����AR�]��)ӳNx(eL[¹$����(OQ>���� 4�$�@@�$z������4O��E)ă9v,�[L��A��4J�Jě�H�[H<�j�2�	1۰=A%fI�e�	�l�2��"��b~
Y9!nfEQ$�g��il��("�	3����a#�Ia��"OT0	�`ADf}���Q�cOf�U�E���I#"������+�3�	4j��_�MQ `6�Ƴ�LC���3~�0�m�4u�&YJ��2q@�J��Չ$��T{��'��Ń�$�^��P
�e˷\K���'j�چӺ-^��'�	��nL9e��{��I�#�RYٙ'�ĐGy��)_�ꉓR�:k`����5^��v �����i*�S�O`�8{�̣y��(a#i3Z4�H��Y��')�D�4%�`Jnј�G9%�B5��b	D�$pL��R���	t�����MU�yf�!����Ip��$�:w�`3�F�
 6A"��c���d�I7ah��dY���!sM�^X�YS1DKE�ayR�.=���'��� ��"���@F�ɶ�60w/?���6�S�O���*@��,M� y�щۂ}O� ��'PT+�ɐ�^����6d[��N>��%lO(�k��]�*��X$g�<>��)���'/��7�Oz�[�]şT#& 0hB�P�!L5e.� �"/D����b�9}y�=Q!��?~T��z&�-?i򢒖|���"|"�D�1Q�܄R1���L��p%M�U�<�",&dV8sGJВ|bt3���j�	{vXc��?On�`dŲjgN�X�	t׌��Of	��䈳C|4�:E�Y]�raI��c��$�'h�����0k��aa�Cϧ5�D�	�D��u[n+-�ه�K�7�p���+!L�B䉾'$d19���5t֕�S$� jsb�j#�5�(�)�'*
H`G�;�z<h3g��nZ����l��rwOEz�"0���	9J3l��=A�ܥ��<����&4Q�jٮ/ȸy#e	@O�<yEMV�'�� `�����I�<�r�Ӭ*����$�B���mE�<�G�3'���P�d5��t^|�<�E �([R�I'*��5�H�2f�Lyg�9HҰ#ū��0ax��g`�
b逝I�
�j冔���>��JM�y,�5���������P�<�|�R���?��X �!�Oj�z��I>7�F��ԇ�g�m��剆.�f�B�	�6�R����<���8G�� �a�`�J�AGh��(�!�V4J�Q�-{nœ�h�hM��$�e�R8�����|���)�矈��ˌS �z��Ǿ>F9n*D��4%��0�\�ba��3����b��<c-E.���� H�G�dL�Y����7��;4 �� *�p>�P���N��!��֖-$~l�QQ�� �5jKy�p�2BGf�� �� �uv�A
7I�3QF�12�*�b���R��*vs�M*	<��J(!��A4�q[Q萢a`�B䉺��ɪ���*�&��72:H���.��q�>��E����)��|{"@X�78�95��ц܁UM6D��х��$���d�=!�8�,�� ��\�%D����'M�iC@�M�li;�(�+R\s�W8.���,	�-`�����C�x�l�ҩ�@.�`2`"O:`�E��/��]����O,���t퉡�zY���S�Z�j�yw��u'���Ӧ^A��B�I�~%p�KY�?�B�(�ݱ*�B�	��"�H0�VYtv$[�AV�Lb�B�)� �%�UjF#F4@e�0�ЈX��=��"O�<cC�%.>�p&"K�>��x�"O��aWŒ�<'|(�v�ظ4V�غ�"O�u8�)�w�J�(Q��[0���"ODB5���@
���b�4�ڤ��"OHP��O-wT~���a�N*V%��"Ox���Z�w�ReoڱC.N���"OB sk��}�<y�$��3zy�U"O�m��`Z9uԒ�c�N�H�4���"O�XJA� �V��-3C,�Qĵ��"O� ��
_�t�C+M�i�V��U"OjEb�k�zo�ِ�E�2J��@��"O���D�(��#aӽ�H��"O�q� �k�9;R'D$4���QF"O�D�ڎYe
�X0憧Pdh���"O��YF�ɹU�R�F�e5��"O�Xa`�AXгl�]'�H3�"O|0i�#�3%��xԍͺ |D�"OT!�/˸K|�(ДJͪ}}X'"O���B;i�
 �iOhb��"Oz���J�5�V����@=mT�ȷ"O\<��N�<YD D�S�X9�=�d"O���b��&���+�]=2��� "O��A��'K�8��A��g��Qb"O����[3-�� ��D�P���"O,WMU�"��4;QE-)�dA�t"O��Ge�@h�dU&`k�1�V"O�8%( �lT�6nƄso<�"OX��cԦB���E,n�ly��"O��a�BX�@��@�A�U<Kю���"O�*�5n���À�Q����"O��y�2 AcW��/����"Oh�:C���!cJ]	dӏ,H�4ї"Od<3�هWDRS*Zd�l@��"OP@�iD!���1�\��"O��#�M��K��w��uˀ"O2�ĩVq�ڙCtj^�4y�aY�"O����=7�P�ۧQ@q�a"O�d������k��K�Y7� 	�"O�њ.S�~by��F�0��kt"O�T����=v�D�BR�*+��9�V"O�M!�L>#�έ+��+�4ԛ�"O��J���h
䙋�i��Xsd�"O9�֬C� ����׳
�E��"O* ��kБ	����Ӣk���'"O�19E�#�h��F��,�:a�""O��K�B��}��DQ$r� ��"O��qŔ�e�X�����$��"Oh��¦1�\�슼=n� ��"O|DJ�+�	D��J�鑥)[^u�"O�!hC=`(���	O/N}��(2"ON���4&�2�@m�E����"OfX�Ƌ��|^�a�]�&F����"O�-
Vn�̾�@��ֵY2�( "Or�3�APN��-�vM�;���u"O
L�pN\��6h0s�U��"O4}�@��Tq#���,��!�"O����?4>�����Me�=p'"Ox�QA���7�J$�v�$"0,1��"O���	ɚv�`UJ��\h.�0v"OV���[�P��A���8�"O� ��C�1�t���oG�G� I9g"OR�z�ʞm�����R�(�1D"O��$U0Loj}A��Z�ɚ@�w�ɓ	��)�W�3� (�����39��3�*ζ]����"O4��厁
?���R����uVh��6�C_���c�|��9�kgo�yK4�=G,�`&N0D�<s��Ģ���*(z�ȃAe��ii��C]��ߓyL�1�����H&��a�֨��I�Jʲ�Ќ_�v�MEk�S��S%E� ,3�O	�y@��Q��0;�y�0����'�"���Dǂbp
<D��k�Z���0���=5� j�mݰ�y��T1gM��9S�Y�-���C�	uP9Kf��0A�6�>�+� �.�*p)���1(�{
��ȓ-�2qB6��.8���Ĺ���w�4m����+3��	�S�{���D��M�`#�/�N��I<Kb�X��(>�bbǝTc���h�K��踲$ͽ�yBDhDF`sF@P�E��1Z�H���'i>�4�2�?9��Fϰ>U؋@�
�Z���b�+D�L�ĄD�r28���zɐ4��F4D�tkq��OV4E�!ȅ>&�(��2D�d���"�p��Bbb\��"D���"�	l>����26�x � 5D��q�牄�Ĕ2��WKR@�B�/D���#M��,����#Y��s6D�`p�Kݞ,��q��\|j�	y�� D���V��#wv^ur�a]1k� �C"�!D���(�S��ȓ�iTO�M{��>D�]�$d �c�Q�u�D<D��jS��'���Cћt4���/D�D�s#��ܬse��<g�!�a,9D��2��c"�P�߳&~�h�d@(D����"�0�&���+�<[�p8��3D����I�F���)S/�(����:D�lQv � ��]�J��`�Z<Ђ
6D��K�Q�]��=B�&ɫ )^`�`L3D��*�C<�Z�x���C�����l1D��i��I�&���i:T��!q�k1D��ذb�)�Sr���Oo�i�r�.6�0y)d�'��,B�X�(}�@�n��*�'�)�̒;`�Z�G����D�U�&I�3�'�ny���\=@d�0���w��J��D֢q�����Ά��')-�<� �i&<��a��K���"J HU�	��呠�'K(�h%g��mIz|�#��7�N�X+O�5�qaI���<*M�lC�c��Qt�D�'�b��@�'��a*�%>Ә������C�ə	@4|r����W˴�gD޷%p���H�d�qOI>j@�l)#AȇL	�́�*�����vD�׼�w���}�e�1��:dt�N�O����ɕ�X��.-q:V5ra\;U�xA˅�_���R#ԑ%Ω[�N
�L�م�~z犂�%��ѡA�����'+��4��X���O���@��`J<�S �:;z�ൢTU.�,A�L4<H��#�Ƌ\)@�%��Q��X�#@�9=s��8c���"�ޅ۷�ʣOȐH�A�<iW��/�*sb�6��X M���
�����F55
�2�l�_V��z�V��!M̆G��0{��'` �Ã<j ��6��-�� z&&0}r��1P��!Ԭ��0�tH��M��4ñXG����lq��жψɨq��L�n�!�Đ�nt mQ6�<j�ǋZ��,���c�PHს��x����1J� qq�%��ݗ&8
�ڴq =�����؈�!^1TULI��I2Wv8�s�|�$��N�v��!��*� � �Ļ���t)��B�j�b��B��`ڌM�x�Gzr!�P 0��A����e��0=� �DD̄:"_�	tR���GW�
��Z$]�6]p ��e@�-xdm����G�a}R�ϲubt�`��|��TAܢ��'��m� .ܟ��������������K���(�4&�L���#ӎ'�B�I;]C�����0p����nb�����\+j�G�t�=c��S�w�LD�&È�yrK�|� ��e�,e~���(x5�Ï{b�|���$]?9^xA�*Їδ���EQ5eq!��'ܦ�;��B�w���!���h�!�Aw���S̈>%��,��mP�*�!��֗J���E�Ӿ3�`�i	�!�� ��pWKI �d%�S��2O�B$��"O�����ʇu4�D����$A"OƔ)��ؑ2HuZ����ZP�"Of\�3$x�&̈́���y�`"OP�J#9�^�S,ԏ>�X��"OY��U<AҊ�£*�D�*���"O4�Z�*ؿ�V�k���-%�,�D"OΩ(F�\�:�ޅJ�㛂8�T+B"O�Yk���."L��W�'s��A"O�����׽HjD����6HƲ���"O\��҅�6&����o���%�эv/qO�uC��{�g�I�-5dSP�H�V�hk���Lr�Cቖ�}ZB�� T���!o�p���&'�|,��	�Z���c��,�X��$�*������O�n%X�����b���1��̰'�6aH��je8C�I��*IX����^����(-�}<���
$
T^��	��8L���2B�Yĉҙ.�!�dF�Jt��M��| �tB�@�8upL��(���&�
c>c�
6ꈇLV���g�E"�h�0�1�"F�I�p
ŃkұsF��2'��S��d��瑽��~b��/YCΐ�S��	=�����0<	"f��<d�eБ�<}R��!E/�;6�O����	����y@;0��9�qY��pu&E ������a*L���)§:�I)BH/;�v�k�D?}����$� ����$n2��³�����k�,"}�':L�����y�/��~`��	J\�+�$cW�Px�Y>���B�� C�0��H�;'n~�x�hZ/U�a2��NK�]���!�Ph)�K¨��<��gF=3A��O�㏽'�>��#��c�BX��"Of��!/�%,��0�%�<�>-C""O�8[5^|���G�B�0��Z�<QCnL�3,Pʄ�\;��(�/�}�<	c��sZ��3AJ�b��4h��[{�<���Z+l���q��~:Y���O~�<yk��l:8���c��4��`0�\u�<qbL�,"��6A\{{������M�<Q�I�O��Aa�	<\�}�h�R�<i�'�oǖA�X��(�K��d�<�AfW� �|i�)��p�[�+�\�<q���+g9\� TNڎj���Qs�<�i�n\�@8a@��p�.�:'f�<	-�[��§���	"T2�@RH�<�5�� �lth�2���seAJ�<��
�fZܹ:�/�<��,P�XG�<9fg�TJ����OPP�l�B�<��F�f��AF=v������f�<� ��������:?��AX`�D`�<��MK+t���x3�5Cx$����gy��M,.����2j�v8SfNPE�"u�K_3]I ���d��zfm֎J�$D�֚TÌ,jW�V�U����vÒ���(6���atOI4,x��Dy�g\uĜ�V��h�O0h%�AI�Y�r� S_#X٦	�'��i6o����u۱��Rv��`hP�e��PzPJX���)��(C�O��]�2i�A^�6� M�A#-D���%�I>Ti�\ᰁ	PΩp� ���b����\�JP�'�\၅�ۊqR�0DLY X�
�dNd e�˺T}d�s��=���7o�%9�R��S!7D��t��O6l�.��%]z�#�� �#� $ѴM�J2"|� �&S�`uI���k�<0QECW�<	Q�D\ڤ3`��o�d���ς�g�y
d��8����O?��B���0@D^O�9"�K&�!�dR�B,��F#��%8�u�����$ն?@���,�0=9vMè/���ԫS7W�y��	AX���TS� êmůKf`0{W�CEh�)�c&��y
� T5�e
��J-�Q��l�(b� ��	T�f�R���cK��0�nT?Ҩ�"��Fl�B�	�.7L2�B�����4��B�ɚ0��@aC�1�lh��VS�B䉬x���ZfՒV-z�I#�PZC�I�=�$�󷋚�5o���E<��B�	�qR8�aP'��k|��af�>i�C䉡qπp1��'JTI�CCX;hk�C�I�9�H�F��XM:��4�6��C�ɯ|�NX V�R�*�QPC-�wN�B䉠o�f*���#)��)8G,D��q@�ƣ	#tmk`̄�Xx=SC8D��j4E2< ���Ã�s�,u�6D���Y:v��c�kR��Pie�+D���%P���зnN�$F}��2D��7�J�Q����荄��uy�%$D� �@[��P��Ζ���lb�%D��� ��/�x0ÀN�Ugr(i--D�����þS<�C���BN�dj�-D�̺�jM1�ԄB�Ή%~�nhA<D���'!���b�1JYH�';D�`�6g��,���0l�ܫC�8D��R�Ô�7��SlV�7��P1��4D�á��q�u��-W&XT�8Q�*$D� I���/?��X�h.QBfl9�l6D�d�Ǫ��<��Xhb��(l�MҦj7D�X���)� �$O)1o����O7D���	��R
�n؆���B4D�0 �N�*rh��QNȪm�7k2D��s�32��������d�����4�s�*���=Z���ie,��|��nԬ�n�z?�DQ�eT������F����/6��m��$�94���F=�u�@��&G�<�#� sE�|�ȓ`�"��I�b$J]�a-������"r��!#�]��9R.и���������*�Ei��J��1s~~(��T��*�pg�d��e�� HZQ��d�O�i[&a#�4ࢣLL�MPp
L21�O�
��)�F6��r�36���H��M=�uitS��q��ʟl�I|n���y��C#�­.���谬�BT౱�Olq�5�e�b�"��0|��1$�ٰ�Y�s�����Ë?�)3`B�� ���<��QHYbN�W�R!B����6L��5!���y�u�� PL#�$|{�li�A�'�d"X�Y `�7��e��'$�b���0|�Q�^���zUK��+������8�*��W��ݱ�+I���ᓦl(^��F��<?�t"%�ۏq����/k���3��RS����:�F��K�'6�vd�1� }�R�'��qrc��`F���\��~jp��
5d+LBȩ�mV���b�bMٲ�,����#5-�+s�I���/*�e;�M�RҠ�:w�|�"V�<�O��'�nR4̓ӅQ�`'|�ȍ}� ��:p�?�'�H)���ޜ6���#b�W��(�	�'�������+���sTHL��<�s	�'"f���%�9���s��&��3�'�� agM�p��rBK�!�j���'�̔H�-��u�(��Q�M�K@iR�'͌}�GH�?!!(� b�R�hbb�9�'3�9p6�K�|�(�qB L>g�Ѕ��'J��j��Z�.P�%s�#�	l��
�'�T��p��=x�bp�Q�ur�� �'j�0��P��!['mۤ�!0�'Y}J���	;�gIBvyB(��',�pi�����a*ȫ���'�@��A?R� -� ��`���Q�'�֔v��K䎱:P��W�h�s�'$`U ���<ѲDc�IE�Nz��	��� D�p�*
r�+�&,	P"O�}��FOA�|�hc��w
�D��"O�a�����uQ��,�W�����"Oh�� ��D�H`c����I�(�e"O�ᓀշxD��K�I��� #�"O,a%J��9 SiF�bs�l�D"O�QJέ2�V���H�g��s�"O.10�a��I��%06�[�dd0�K6"Oޱ1�VۄE2�d�k�J�d"OdQk�Z5Z|h��ݸ�6M�"O|YJ�	M<n"i���@~ՠ$�"OV�(R��������H���Ҥ"O^��FμRHirS��wd4E��"Oxe�o]�0�LQ�T���m\f,�d"O~�1W0E���9f�Ҡ]M�\Qu"Oq[�"�Լ�V�O)d�N�&"O�qr��-�]P�,֥,�	d"O�1yW+�q��Ѐ@�������"O4���Қ}�����=3�@m˄"O4�XbgI�14�sB�ϸd�f�c�"OF���$y2�b5�˻i��)hu"O>irtϓ ��(��ќ	�L}��"O<E:S��}��p����`�X�"O�x��D�{�pc��
a~�4R�"O�L!A�?'>~T�E�>i�`(u"O*�9��3Ll �Q��n��t��"O�t��/���2Fؿ��AJW"O��Ǖ�f��I�bJ3p� i
�"O����܎9��]��N�����B"O"�@��-~��
uͻ.�`�"O�j�f�R�^�7n
-q*��"O�%���ݒ�(b�	�!���"Oh̫��O�d>������J��(p"O����̔7�\��#ӶJ����"O�X8Rc��=<��C�g�	�ƅ �"O��t��!G)p��g��֮5��"O��R`�:࠙��f��hc4�RA"O��[�ک,8A����6 # "O�ؑ�/�Rh���%��)�	�F"O8�A4�d0Ё�p�� !�z�p5"O�A)S�"x_�E��#֧�q�w"Oĩ�� ��1��T������"OD�a���)�њ��Y���|��"OƑ��],?X����>��+�"O"��E�_��"����?,�h��W"O$L
uCA@��d[U�<��t�q"O�4��K�"R��@�LǱ}��i� "O�q���$g`�(�7b�"�v�`s"O ���N_% V��*�ª&��IR"O�H
Po�-N���۬w�.@��"O���PL�4A�d��u�T����{�"O���Ɏ�Mᒴ3��
[�`�"O�����i��r�5[�	@�"ODٻ��%w!|�*�k^�$P�9��"OD]s�d�!�h�:d��.@<�I�"O�ա+7��(�[=fA�g"Ot����\����ô:��"O0a�r�	�'ˀ��P0t��"@"OX�1�$�'kgԋg+M�<J�"O��{�A�$x�y�4��$��}��"O�)SU��,dA�p(�Uɼ��""OhX�&`���A�:XbE��"O������gS�L��D��?�Z�s�"O`9�v�/k�qTi:|�J-�S"O� �㴌�*u����	�|T�W"ON��7�� 	�Q����	�h�A�"O�K�Oݼ}�-c(ތfD�t "OP�"ť(��c��<P3"Oz�"2H�)R$�AQ��%,
ઠ"O�2'ɬ\Ė-Xe�=RY �"Ol�Kb�˞��ї�ʺ'�,}�q"OL�%�%2��mqU��|U�"O�Pr��R���$�m0��|qP"O���#+�
<P��,��-�v��T"O�
E��i�V��r엍Y��K�"O �1ꘝG*u�ת�Y�X}*��'pd�.OT�����*K�p�5k�m<T�"OL(�W�p�v�Ya��Y���_�ODt�ٔ�ë���j�yE.��'����ЗY�b9u�n@�(r�'�\�%E���D����5c��)��'D8�cH�	��Zc �5UT��p�'s�h#��/e��HY�K�����O%��	�@��aB��P��
\����	O�/��*�K�"
Ъ��r� r�<!�*��N&sÞ!��,p"kd�<IS��O,���q�ŉ�k�u���O�������|�0�#��3b�Z��'y�C����R_>Z�셪�'����DV�_�����O�D���'p�5CW'ׁ|�J���)�`���'��I��-T��P��3Ӛ����'�*�l�D�,sf��*5[�u��'X4)�G�Hz�)֠B�\X�, �'��@�G�5s_`��f��&NX�a��'����*�}�]�1��\��5<O~���H� F>f9Z�e`Iҷ"O��Y��&�P�$�f].th�"O��叛$=^����E�Y��h �"O�u����7�\����:' ���"O���e�??P�ȑ�9Tu��`"Or1��䟺�dPqMU&&g,�[B"O�1�th�5Z��ٛ&y^Αx$"ORA�r��`�ɓ�.KXO�p�s"O` ����uԈ�3�TF�$�"O&8Ǌ�D{V�@�ҏ!�̕�"O,�c�灩x.LicMQn�JQD"O�b��D��X��3�T4O�̱�"Od�KT��ܬ�D��쑁�"Ob��qJ�$UN���φ:
�(<G"O��r��Z
Ȋ� Ж[�N}�V"O���@��s2�k桚+s�֘*G"O����ɕ7��a��j�clM�"O��b�@�>I��)딊	�kMrY�"OșQ6k�{䱈��	K�x�"Ot�x&�]&]ي9	��5gpM�"OΨȷiD�+P8tRgbˇxg��(V"Oa@S%҇}�Pݙ�]���e"OZt�����K�*.���u"O�Q�����
Wn�)`�Q�2"O�8Rֆԉ]�Ԕ� �H:��m�g"O�ls��>�t� �T;Q�
��`"O4�K�ꊭ��4
�5rtZ��3"O"�C�)��y3 �C�Nv���"O� �AкxbpQ�!wm~��v"O�a�`�#s��Q�!�)l�Dp%"O��k���12��e��ԓe��Rv"O�H�c�k~ѪpG�/�"O� �5�Ђ??�2�{R6l�v���"Ob$���3
\P� �j�8(0"O��jU�^<T� �NH���ث�"O<tR�M�:u^H2Í�1$r�A"O� �dg�|���G�6
���ö"O�L�?e@��l��Bdr���"O�9�4��T����(�"k�n}��"O %�G��cG��F\ �"O��J�[�5 S��j����"O�e�W`R%E��9a�k��Ll8�j4"O.��w�xx[��I�Pl��"O|�3ᄊ��(]MA�'�Ԙp"O�i��ȯB��"M]G*��"OBL�� �I�\epS��R5:��"O>	ȥł�5}"�S\t"O8�Zt D�7e> s�̓���� �"OPȹ1�ks>���Kɫv�H,�""O��wmX�:@��G�A�s�X�r�"O��Sec�I{����ƹH�- 6"O���D;"U:�ƁB2"�H�"O�i�U`�SHj}�􀀽p�|�V"Ob��UcN���(A�/�5ҷ"O������FAAѢlFm:�"O�}q0`	3�|��e����#7"O�|y�E�@DN���kU�S��<��"O>�@��P�aJ5C�	B�Jl�%"Or�pv�_�D�h`�� t "O�`@�D��ou�Ja"Bxj� ��"O8�
��϶.��E���U�,�
���"O���F�/��F-�����"Oҍ����<C�{���z4�X�q"Oh�@�d��R�T��1�N� 株�"O�q+0���8�����h }k�"O��2�Ɩz�cs�*"�D��"O����G?Wcd�+���=]���c�"O�Ih	<tƜ$"�D	g�D�d"OT�3' ��]�MY��	6�j���"O:��-����W�n���U"O�I�iӤc}V��G�MИȺ�"O\�Ɂ�{��`�q�Z�[�`��@"O�Y��_����5���r�%"O�q9��PeU�CT,�L�0,�3"O�8۲A\�m������u�N��"Oh��(bֈ!�E�$�V�h�"O��s&��<yA���d֘6w2��"O� �ª�lU��6�Zf>�1�"O X�4��=����A6 �S�"O��iSiL<E�%83D4p�t�"O���Rぶ"h�x8t�(��aS"O�!@͑j^��A5 ծ�	�"O���mI��dB��Dʆ!J�"O����MJ���|+3�R8_��͓R"Of�'��8��E*g�ƿn�����"O����Ƙ�񐌙�&��|�TY�g"O�<6I�<��!D$H�@`"O*��N��;��\���'Fx���"O�ڠ��)D~$
�k�
)����"O���kZς�@̏:��([�"O��q�^�n���c�	Y�%R�"O:�q� 
  �   �	  �  }  8"  
+   �pA���D���\�'ll\�0BLz+�X @��e�2b� ��/?~��'��̘��BF��	��Wy�(C&��_�hHiW�'���"fՎ>!�$ѕ�/��a�7�7t���'	�j���W��i�ȉ21�Q`���?���䓫?���'�`)�@,�yJ�Ӂ� &GD��ߓU�'[�Nɣ"m&H��(p� dX�{�:(R��B�����.�C�G+S���SR[�lT�'X h�D�	�'�n�SK~z��ޝ� ��%�ǂ&R K��P�<��$y��q��́ ,ʡ���a����?�,`��Dj��C�Ur��a�<��LS!~)#�bX�
������]�TQ���'�$��>۰�8�$?l$Q��D�6<�}�<��?}�@�Y�\��ts����-�1�̋i̓$��1�0�3�D�83�da�X�x���(G�����ȓ���A��Z�"L�T�m��'K5�	b���On�U����?e@��O����'�d<�v�şjD��B:~\��i1�Iv���!�ɝmO&�i�4,�H�"e�\�\��T95n��<Y�i�X�O6�R�Y�
�	H�`� `� �Th}���C�Z�uaL�{��S�ҙ,H��ȓ)��a���6� �+B�Y�^�Gxb�'�
�)��J:R���Iw!ȁg�bx�'ia�N<h4`�(M�d~؁c��Ad�	��HO�i&�$˥��E��8���$A����iJ�e�hX�R��?����?���4C2�á�?i�e���0��x�����B�2�&OD��r<�U��w8����\!:����2X�B:#���͹v�W�D�@��5IJ;]���D�5(��8cL�M9���ơ��M� �O`�D�Ԧ}�	{y"�'ȱO��p�F+ٶ�
"iN�.�r���>Q���U�I[�j�����<t�����1!0�M>��H��6�S���i��EdF����䳴�_'z���Ь�+\�� #�>�&!X�W!R��4X�&y�K~*$	Gފ��V�S��1��^X��T�<6N�'r�K�dA 3��M�oЎBR6�� d.l�I쟤�'�y �ǅ	(�~��� 5j���'-��'�O��KF�\_���.�5~��Y�@��_���ɀ�H� �)CV F�b�I�kŅ�z�Ӕ,�O`�1���.ڋ7�48�|�E*Z��Q��$8Ȑ��D��)5DZ$�g��Y��޸bBZ�0OA}ܧ�������(چ4��If
s\f�'�x��� �S�'2��`�M�J�Uh��S	$�,����O���8�)9��قz��aX3E��P>Ń�@"�(O>��d�M�*����[�w�D�G/�R"=I�O�Y��a��nh�XH��4Y�`:��ӮJub}����O��D�O�����űP���d�O���O\X�GM&���J��ɛ_���QR>�ػ�ē6W�P<��M���Q��k�5:"������&Icb���0RE�K�Y�x8SN(t�AnD;l%�ȣ�H���OB\X�֬d�]@f�g�A��\(j��@�h�ac���'� %�O�b�'���'D�F��*9������eľ�Ѓ_Ĉ�?���`�i�`�R@�
t0�:�!��kf:E��2�yb�L,�y�I�����N�Y��~j�!D	�4��@��4���:����6��г�.��t��O X)���3���<�6b�:���Q s��@M�@<)�$�'/KZ-Y��j��x��Ր*`z���,O�tpT���k�<�Q��D���@��<�	��6��=�D,�4l �6 ?Zb����	��QT��9#,�6<�⼂�˞�*���=��/��^��1�`��<�ش�*h�X�
�}x5�ֳd��u�!�'/���8)�>�I��'��,9+��J���y"�i��9Ђ#! '�5(FK�M/�`j	�`!��Bs�R�����G��O��I�σ���\ZqL�.�Ju��'��#��?�R�in�&�۾��ȉ�`ծq��	d.��}B���?���O��':��cC+�ZM�q��\�r�k���9�S�TC�
��� 
�/Լ!^?/>����'{�	�"E䐦d���4�	Q��J�$kכ���8\i;��Q�P&�I��@�`�����O:V�X�r��{��O��'�F�C`�۽S�N�+T!D5hf��O<�E�Q���O<|Ի0d��)��D����hƈ�L<�$��Ο0������	Q�'{v�Y�`�h��	�
�l�PQ�=��ǰ<��ș�f��pf �5.������HO�?YT�JT䖬3��4+u�E�:&D+T��OD|�͓�?���2������?Y���?���*:� <8��a�=|����$ �)_���a�'�,-��'�@�͋�G6��D{B�Ȁ^;�\( X z�*�@f�Hg`�y��>�4gA0X����'@VEZ�,�:�Z�+�Ʉ�/"�d�O���O@���)�Oq��I�Y �*ɱ-��My%�L+&hpР���xrd�28"�MpE,��Hij�Č*�?�%:O���C����T�'�In1,L���U�&��⮞�<�j�(�"B����+���?I���?�WG��T{�������T�L�zY��ᇶI�����J\�Z�d�	D&^<r:��"���x�B�ʬC��2��ԸO�pQx����v� ���w���#�L>3ʖ��FR��d��ޣw���B˦1�4�?�/O6��<�	 v脚eǀviֵ�$�-����q�'CҴ@��$M��� g�)P����k�nr��'"|���Q����4�MK4�ݨ2K0q�-�YrN��2E·D���'.��'��^R;�������%+�,O���&T��P:�N�e�P�kT�'� M�'���+�~�!&��:0J�:tk��ayc�,�?�e�i�6o��U;QE�y����Ai��|�ŉ^wy��'�O��z�n �q��I��H�����Z}���i�1����� ��X'��hS�A(u0O\˓7�1��D��?���iSx�6ɉb����-�ں��W����R��I��P�j�3|X����DW~��]�T��"�?թaCJ9L`���UƗ3�*�Ƞ�#��2,���FSB�?�K��h�8�Å�<����3��K�ix"�yӮqo�����~Z�fMZZv�;VN-m6����d��?A˓]@,pg��<&A$�R�o��4�S���?傑!1�I��DA��@�W�ݩ��.a*���ו�?���?��O�:{��OR���Od��߂W���[ů��>1�E��..L����=)��tH�P� E�L �=�m����h�!s����`��G���yK��������/�����.y�B��g�2]r���'W��'v��P�����v��s(ڗ~���1E&�e��5�1�]vH<��K &�ġa���	@��:Q̔谚'%0����y��������Gڰ���&E�m��l]�M����=���i��d��J�0���|��1}�NQ/D�6�DE!-��y�ƏJ|�X��ӈ1��Y�EIU>�y�FûrFU"�
��+����Ag��$�u(��rH"(���0�{��?��LY�4 r��eA�=#w��.Wx�O��GzҤB�(�6�D�^�e��lŏ6Ɔ�Z��V��6P�����J̓d|nh$?��P+�!Xc�i����PQf��!�4D�4s�j�(,�Y�p�Q:
���3LO���i�NL1Txѓ!�P�)�x+� 1D�d� &� L�Hk��
2�h� #����HO��J$&h�Cȁ/$8�+b�3"�.E��ϭm�J9�<��)��?I�T;��2��Y�l�չG�Dk̓sg����2�3�d�&%�e#�c�t\!"Ի2}!�$��E*Q�%D�(��3���#H1Oj�=�|�TH�Zʠ;�/A;+á�	N�<��-إF�0�+�^1�� /
��HO4ʧ��O,���*�(X�#�_�`�[2�'�Tpy"�/�	�=�d"|b��0w��I�ӭR�L�b d��
�v@s�H�d���:� ؄n���R>#�rH��E1D�4�D�y��尲��i�f��0���<�������5gX'ڰ�qS�^R�<F��n���ιXt:1PgB���s�O0Gzrn;����1��($�)O�x�Q-��8���D�S춄I��B��	v�|"bQ��a���<�,y�eH\&�yRL/��%˂08Z�Z�œ&�ybJ� ��� `M''�x(5H�J���/����"�<^d,B���.%��{b$�D �h��3��"nFeIZ Z��OH�Fzr���%r��ą��!�sn�3W��Z�".��E�8�3��Ji̓$*��'?��GgU�[Q4���ƫ2���ɳ�.D��ӷˈ=�2�b3�D<|���v�.LO��`(2g]��ֵ�c�A��UQ��'D�t�G����m�  ���/]�P$Z��Q���?u#��P�3A(4�&L�w��H�6��?�HO�u2�Gf̓Hh]�/�`�2�kV]fl���2zi4�<P�	z���>�O� ��X��&d�P	2��=�� !�"Onq�iL����4�MRF��%�ŞHc�C�3 ���#�	�~5�ȓn�a7CKm��h)��@3F��y��$�|Ұ�dF%k=�%ap)�;��8C����{��펭yh�b���S�(�'/t�Uq��"f����� �`��JZ;g����I>/�T@S��ݐk޸"���)_�B�I#����@J�>|��$z �҇sK"<�ϓx�
���m�hͮ���@7"L�ȓ9jn\a ۨhb� c[2�ʭ�	+����K�'C��O����*�8q$�h�J�Iڹ��OT��3A�4(51O�IBB�q�'��]�E�]4^��	����A`�'|<�&'Ȃgd�@��C��>��'� Dy�dde;��^/����B,�Uh<�eV�)O,����_=]���#�Q~��\H>�·�FX�C,�8_�Pq�1%�x��##��P���T�?�bDV�R�ĭĬ_�A:���sI�v�Z�u�t���D�::�OH�@7Ļ{��TP©��eÌP�'Z���0�J�3,i���=dP�	���'� )P,K�L�� �p��	A ��	�'C�;e�g�T�H�(*V�D{�re/�S�/0e9|T��N&m<L���8vMN#=	R�Gc�1Op	
��O��2f.�??nh�f���v�����!v����L>�"�ь+p�}3�ǜ/�~���I�<)��Rr���3 /.?���P��hO1�v�a�E4se���)�[����P"O�͠3�-P��8y&,�&�)�m1����k�3����	e �JA��J��Iv�`��y��\���\H�C�P��Qcʖ�V�JY#ko08B�'�N=C1AN�-�	�c�+یM��'T��yEB։PP	#��F� �(r���+<O�$�c�Q?S0��BLI�N>��"O���F)E�Eu*l12,ϬT:�T03�'��4����J>a��<C��d�ܼ��mؑ��g?�a��l��<Q��l��m$�p�*ŭ^�4����T�g[���r�2D���cK�_���A�ȏO;�,Xv�"D� ��
�A�)��k�}�\�0�SZh<9�*���et��_ZR�i�HJg��<JI>3G�;�00 ��yXH���� n��bt��`�ߑ�?)է}�ȹ*�eF18�"���q�ĉ�B����P7�O쥊��S�Y��G��Z���' ���j�/fD&���S��d�ӓ��'�~�t 
�j���ȓ�� ,�'(`����&��Qz �S0g�B�3�BH3�S��ϊ'L�Č�+do�anJ ���!j�f��<���f>Y�a���r��0Bҙ�Xq����|�1��t��/7�3����\��PQ�d�Nw�8+�͝:
!�dǄx� �asK&@���R�D���1OR�=�|��B��l
���sM�!**�9��?T�`Ԥ�.FH� b���+=����f�'8哶��'JX�قOŨe���
�'D#��)��e�q���#�>����Jx����k��#�Dj6�B�e1�QC7�Ov��.��t\��`^03��#"O��"����!��7 h���t�Vx���eP���@P���ykŀ:D�8�j��k������� ��IT�O��'�x#=�1�|�+�n�L)�C��m��	�&�(�~rF�u�� �yR��ݦM8�|B���U��|�3*N#���K����y2G�Anmaf�Mi�d;�,���yBJ[3. �1��//~B5��ʂ?+:��䇆F:�h�&��a��w,95�{b<��S81�v��5`�,CF�8�@'�9�O6�=��X���U�3���g�X�:���b�]|�{v�t����x�^�`�%?�ģZ?Sw�������q�H;sh/D�� �U��)�b`�� 
�T�6��#�'�O
h�耕+7�5�X4��"O*b�C_�*�0<�E&�y��y�a�D�G���)ݤ&Q�<@��\K"��\�HFz2"�2|l�c�8���2M{�f�*[����G��(���3�6�I�`W8�	���|"�6|�"��	4Nv�1�Z��yE �1`BM�h�
��X)Ao��'Mўb>9�0��l��-���J ���,D����M.n������6H0�`J\�' ��1��'%z�C�b��8����I���n�HK�B��>��7 D2\��ŜaW¸�o�+X}��e�9�OZ���-[�7_�|r'o��.�8w"O�<�'��z���`M�}P��0�Nx���O�U�jQx�d�/�8�@`�:D���J�b|d���DW�m�ԃ�Op4�'��"=�!�|��?NY��`�7b�R,"Q�
��~2�M�cB옉y��O
�K>�G��B��㷫�J5��!n�m�<�uƆ?G�<�@aC�=TTXh&�OR�<Y#�A�kf��2iO0Ĥ�PD���x2ڌ!���0#��$־e�'����=�ǝ|R
^1ͬݹ �"��,Ki���'? #=��W�\Z�l�z���â>\�@* ��䓣MVc:�	9X= ���M@���|���c���c�>�b�"OH�k�� n��ѕ�$�B�'��OL����>t��5�scԮ~8�	�"O{��%?ۨ0��V5z6�x���Z���ɞ�Ud�2E#� �"��C�D�Σ=�Bʞ�f@1O��B�O~�b�@�=c���rlA�%�����d˺pɉ�L>���0`Ȫ�����&n�8ѻ���F�<��.�B�A°��	m 	'�E��hO1���򗩂]β{�&��p���1w"O�b��ؗ-aڠWG� w�E��j1����WR���^�ɖdR^�h`��
S8���l���ڊy"�O%��F��D˝�(�\���Y>q� M��傩c��Q��'?�5{$�ϼ-զE�v�T�m*h��'�$��GE�c�������d�0Ƀ��4<O�ŢtNEb��@*��z��1�#"OD�P��N�KS�x��H�U�XJ�'�p�|`����L>AF��P�B�A�V�\���a?�����=�I�>��="��%�Xc�Dج*Y4I�!�-R��1D��R&��:�&��*ōEN�ҶB.D�b�E ~����ADB�B�#g/�ph<����/����ą+�T8��[��4;M>A �ȟ-n( [�G����B_|�������D����?�����l8��4�:+��|C@�Xt�I�
�|�Q��ą2e�O�bTHS��&_̨�:pO�ap��
�'\�R���>h|�����pBn����'S��CqGL^<�so�i�Bȩ�'6����㒜L�<4h�O��a��{�R�,�S�Ĭ��zl8gCˋEM|��
I7l	ў�+�_��'�ȵϧcb���S¨B\d���D!d�Xhy҅B(����}&��H��]/PŊD��dKa�� D��H�K�sѨ�y�L����4�	l���O�`��u��Qr����dW$,�-q�'���Re�Z5rZ�����"$�qp��IH�t5�IqP�Iq��W�^���ǅ�Un�䖔h��(�<)��6��<��L�"?�M�U�H�7\B���CP�Z�^���+d�%!�B�1X!e� n��L��B�I�Pv؅hׄSo�KK^3d*�#<��F�r�; ;\Xj�d·��+ D� Q��зC0H!�ˑX��`s��O�u�'��#=q�y��T$V��D��.u�Uc�͞�~�̓�-"ΉR�y�c݉�!0��N���b&e��P�֍�'b�*[H!�O-9�*a�Ӏ	r�� 3d�#0!�� (0��!�+�Nm�BF�!Ou�1�44�IWjmK^�E�D�B�8��"|OT�%���.O�E�$�"� �z|5���%�I��u7�R4�?9�X�?F����>m����R�m�V��c����)���F�����R�90�<"E�2�!�D�1{%���!�(�u᧍իW�az��D��ݸ!l�r� Q�W�B�;�!�$.C3��PŤY;aUV��$
��O�	Fzʟ��G��3S��\�R`��q�j���?ړ$i,��d֙��TdB$;����h�����
�g�1OL)" �)����h�tzFX�V�����K�{x�5�ȓaȆ���o��'~r)�%I��(�<���逴�<���-&}�E0��J�@!�ns���#��N��J �$s�X"=)(�d4�?ׂ=p��j�O;v$�H�P+H
F/ʔ���?9�<����W�i`��'D�V�+1�;�l}H��\�	� �A芄%�z���>A��	�u9d��ԁ6�L<�ҧ�#ej��c,�9y�x(����<��:�� g}¦���Rb?O���Ar)�!�B�G;\��͛�&	��|�'������|Z��dsAجb�ڪ}��(��4�!�9��I����$���:`��|��%|��97�6��?պ����ďKf� �+D�0��@�� ��4�����M���?�����
%�
�$v>��@�Re !q4e�
"f̬��L[ ��!E�W�Aad��H��x�bY��ն�̻`����rĴGQ�d���8�$
W��G��
�'� Qɖ/Z��Y;6dFWjV��A�<��hO�b�B�f�ON�LCa�)A"�X� |O�%���@���f$���f��='�tA�*?�	!l�$��Ry�J��매M3#��$}�ypHPs��W��ڙ������]2�Dk>ɊcG_�8� �:���@F.��7�2l���DI�����#&�wb�x"�Ɏb�l�ul
	b	��V�W�~d���G�RA��8bP�����O��('Z�g	�~bR]A��\���=a	�sR��95��U�x������9�?W�~j%J�ِ��+i�$P�qN@j�T����u�D��OP�_>��ٴ�M��1hӰ5y4��a��H��,q�2�'���Ō@�>O�y�˖i}��Rk�u���?�C�O\	��SLDp���`t�&�R����0.�R�$F��. �?�`�A���z���zA�E��ē�����ǟ�D�t�i"��p �|EV�!�ɒ�<�X3�'����a� 5��y�@%ռ3{����]"�OT��[Hp �
��R�R�'� �t��2Q�,#��'8Bޘ[��7���>�D�O(�1[2P۰$^!)p�#QhՉ
�|bQ�@. ���!�O�!	s-
:Z��HN?O��+d���E)&�@h��.AN�r�*��qf��PWD���?i�bڳ@±��'���C1E�R�*��ԩ�X���#�h�O4��"!�i>�Dzr�»vڪ5!ŉ�4Rt蛔�ϼ�y�� =f�m8cl�6m���#)���?!R5O��2���!�IT}�#ב.���".��h��Y?p=�g�ۦ��	ݟ���Qy��d�8��8▃Z�*�n�[1�ܐ��,q1��TPv�-732����:v��`R��9RVuk6m�'�d��N�=2� 	"tE�,ְ=�w�I@��#ӳ<�BȹU�N�;�$i�	��G{��d�?��a�/�����P��M1H��{�b/�䕙d'���a������%�L�qO���O����&3��ɇ�?�<�푬Q^�	�uG�G��O`��y2����'�r���Nٮ9d,�6�Z�⌅�:�����k��H��C�$�
$��I@�U�*�ꆧD�C`ꡒv摋t��i��b�=b3lM�hK� #��N���?!w�)�G��q� b��4RuP,�t̕��hO��A,�c̓a��S%��ThP�/�=��jL%e��<���9`��>�O�e��� V��XB����G�D��"O��@���J6&lȆ�Ňv��m��(�S�'+�� q@���-v\�7��I���ȓf�Z��)a4�!ZJrp�ҁm�'W�S���'�|�@ҩ�^��a�'1�1�'�����?v   �   ��@��?d!�$�ZCE�ԬG�Y"�k���=9L!�ĝ^ҪP�N�;^\Ppg	�V�!�$�s�,��ӪS�k�Mz��F7z�!���E�H����*%��,c'�W�GT!�D6�Hс�IP��NT� �?FH!�ѡ>yLyⶅ�W�X�{Pf�h�!�d�i���r��%R�b\B��>�!�d�<9j�p���2yv�C�~W!�D�1�,�r0��8ZZL�j�F�
N!��[�p�* (ÉX+�!��!��V+g��^���o��FL�ȓO��h:�J/�ܽ������ �ȓJ�����pg�)��U~�L���S�? ��2���D͖����~�:i�"Od(���6 ��@�f�O8�؁��"O���W��-o�P�D���N��"O�6��M� �%x!�!h�i?�y�K=_�j���D�j;���.C!���4o�F��a)�*�,ˇ��o8!�$@�!�`��T�C +��E"4@��!�D�(��j#GFE�h�0�o ��!�cHP Q�ь"p��8�NחXA!�D�S����ݑ80��3A'�f2!�dI5~��y5J��q����^0t!�WF"��D������7E��T!����h����+e��$��$�!�dԵ>�� K0�$X�Tȍ�R�!��W7@Sm
�*��@F="�!��R�3r��8���W�.��p\;�!�DP:	�TB�g��*��c�4j]!�@�JXl-�t�6�.�{@���!�d�gU05+�к��Y)Q� #!�d�Coxu:p-�j(z�n^�+!�$�1I���H�^���I&�� ^�!�$KS#��Yu�[�>�d_:�!򤈕+uj��W�6M4�\Z�흃Z�!�d�%Q| ��D�GD�+�{�!�]�0�pg���\BuX3!�zH��Ռ�.Z8��&`!�Z� $�q�7_����,�m!��[�'�"d3��&# �C@�$H�!�D��t�٠R�9�JXc���!��&G� ,�Eцk���z@-�!�d��r��"�?B��b�� Ff!�d\!1�z��7�.��g`9B!�D�=�f�S@���n�.V/!�D�iP%��`�>!V�� %���Q�!�dL7���x�
[����ω�!�D��^�����!	�*8CT���!�D��.Q8XyvK�-p�╺Ӭ1!�dZ�;q^!� m�e�8�v��!�8E�H����L)h�X6�MQ�!����		��Vuan)3�Fܒ3�!�H�|�� ��pW�I@1�K;X!��P�2�YR�ܷ~U�1c�S�4�!�$X<1��	�᭜�?aJ�ʷd��!���$4�!���Q}��e
@ !��xrx�`�+F�+J��cʭ�!�D�W�d+6#K�:��r�I#t�!���G�Ȑ��P�u�ԝ9v W=:�!��ߜ$jűT����8D��%�!�æY.,��̔ 4���I�E !�d=n�D챖I�$6Dj�´��<'!�$m{�e�tn��'�:���Ў]!�$H����I�`y�HJ�L�?�!�dM�g�L���	c�ī��3�!�޺��h�D���B�|�K��V+\�!�$�	fJ�C����P�.�Q��:b�!�@U�~��Ba�?g(X-ɶ�N�w5!��t�� R>F2U����	*!�dG)
�T��	I3/Y�,���U�G�!�ć���\��4-:6,H� K<l�!�d�g�v�h���f��Y��\)6!���?s$`�*:&Jp����N+!��^+8!"dh�Ƭ8B.��1!�K�Y��8s�.]�:q�6 �	7�!򤜠v"�����Q��
���Mz;!�� ��34k�'���RE�@�Ơt"O�i +L�4e��n�w�=�U"O�ѣ�I(vi�@R���X�P�!B"Ont����^�Ƞ��I�C��5+"O��(R�O;\nY�Q��5��\�G"O��32��>I ,��Eg�������"OJY
��D��40���_�N�v�8B"O5�6�� "3t��'�=&��Mxa"O`@;��Mt��煊�v� ��"O �K�K�	R�:�$\� uԌq�"O��ȵ���p�;���:t�"O6D�á�1V,0�G��X�V�#�"O�c��I7l�m�!$� &;�D�"O6uS��.��[��]���3�"O�e��ѥ_Jt��3��6E��;U"OH�(��)K��¢��-&@,9r"Oj�Z��y-R`a�	48$�|J�"O����y�R�:Q�ާX �-�`"O��G��8e���P)E�e>ɚa"O�4{��O�!r�!!$g��`���+�"O�)H���>�\ G�s�nq2F"O�Eh�J�W�䁱$Բ�@��"O���Ak�
?�|#փ�}2�Q��"OFP��ׁ �vYɆ"T�<$&��"O"�8")�)�H��A�A<`�P�"O�a�⅍ t��6��0N�@)��"O��ѱ�USƱhr��T��Ժ1"OzX�C,�Y��9c�O"Mj��96"O�lP��R#�]��)�SɶAs�"O�jfƂ[ufEk@Z�}��4ۥ"O(���F֍[��%3@�e�ZE�f"O�CQ�\/R�i�Qo�9\�Rpb�"O
�ޚ&�Yk�,�Y�jM�c"O�q� iFq͠ �J̸v�L�۠"OL�rt��/�Ni��⊪J'Lے"Ov����u���a؇-���xvd[A}��'���� #G�D|�Uo}�Ʃ��=S�+KF;Y2n���?�C$��=���4)ˀ:�l�0Բ0�7o<���G"��gC�C����'x����k�vӚq࠘8h|H�Q��y�I@��?q�4���O��D䟤7�[|J䱋š�/sG��FL�^f��D���Y�"
�(�R$[V�L�DМ,����CN��MKN>����/O��pU���Bڞ��V⛯W�2m�͐ ��mS�'�6���?9�E�[N��c�tL���FIg�RP4�ĠFK�}-	�V$J�)���T����&lK5m\H�h
�I1�h V�1h�n�rU�ɨt��7��kR��1��Q4E�I�&CJ	W�P�	��M����D�O<��)T.P�dTL�9'v>���a/9���(O�D�?AUN�yc�Ij$�1�8��P���4br5lTy��H4�P����
a��(���ʴ\����[);$�'����?I	�b����o�,y'�P:u��@��21��K�'��uJ2"�!�,)!��I���QN��FtcL&T~,���%�V����D��[ "�'�7M�O�֝�fG�9��f�fA��!$�)>@������'}�)�'p�t�
s*C/qER���'	<K$ƴ&���������N��7�<Y4N8j`,ϥy��Hyd9{1����M��@� �z 9����6lZy}2/�{+|��1'V�o�"q�o�	�@��G+���,��lt�?�JsMQ���;zn��B�"�	Q��$mO��4ҕ!IL�e���B!�=4Y����	�n�&�M��%Tr]!�͑�v��	�m�$�$�O�oZџ,F��D:�����V&���haM'��Ꟑ�?y�}�50����tJ
/.\䫔!����'�ɢc7��B�4���?yK7��UfT��֣C}�܉��鹟X�'����4g}��#>QԭD�U���CsE\�9��Z�b�'<�v�	��� ��Է/��� �+�0s��:	, Ȅ�F�	2�F+� ״5p$3Q��b�X�h�h�s��2�S��4I�d!΄Fx��%O�,�:eZ�4�?� �H��?��S�Y�0�I�s��ՕK"Bi���J=>K�m��f�1�hO?7�{s򥁍�`X�%ڠ�\ΓXH����i��'\���?e�'?H� �Ͱ�ՠ ��ݪP��i�J��Ub[�M+��
��y��'��A��Ee�H�S��
V��Dۧ�P9qlJ`p�ܡCJ���n���t'Tg��x0� ǣR��D� JԖ]6�q��M��S��'����4a_�(r��x�6l�LL�S�v�':O��$�OH�O��'2�Kڞg7���RnީŌA�Ǣ!<O���?��&)h6���ү��,����/�x�d��_Y��d8�$y�pX�I~}r�E? d  ��ڑ�
oqL��R��+NE�I՟�����M�Oq�6=�$t�A(T���R��'L���ۧL�O���-(I���, �x`Yv�'���\T����j�%8�D���lD#�N�{��Q`��PZ�'�B�ȵ�����Y�����Ĉ���R������X��q��F!.�X���U�*�����?���?a/O��ȔoO<P���O��� (,�4UСȅ�k�Ə�5F�L:�������O���0���Y�G��,:� �.U�����tmj� E�2r?�� �L�p��]I�-:�'l��L b���*��T�'{�L�A�Qerj(���
럀�	ߟ���m_�t-�8'?������33���l��V��(�$k��	����� �4����٦��	���Ӽ�I:!)��7���!�^/�����I��?Qs3?x���)IY\��43@11m~݁�S�W/�,�%�K�4���«�?4��z�\����g|| ۴7A�'��OO@�{�l�5wwX��� I�_��U���Z���vi[U�����ޟ<��7�M�,O|�1G�T�8��@�$��YZ��`}��'�B͒�~b��g`vd�O�Ei3B_��j��1zztQA$�6V��7���y�'�;7h%�	�"`@*O��ɕ��鱄��lfx����;N$LuA%Ś�@���ԟ �Iğ��_yb�U�L�t�'�$4�,T��td^�qc�X��'��6��O�B5��C�O~�d�O�I`0�O�@� ���<aU�LB��?+x��`�0jR�z�4O��2` ;�u�@͙~X�u�O����Q[��r�eS�K�^l��"�"t�����Nm�p���Ο���?5a7��c�s�I�Vő�E���w�r��eʃoVğ$��ϟ8@$�&�Mϧ�?Ѡ�i�j�/�y"F[��lx�׫�_�z!���r`����'T4�
�!ňd���Om���/"����'d��A�
�4!��V��N�d������	�{�z�*O��	Y�%n��?����?���1[Z��cGŊT}z@0D���?�����Ƀ%�\��F��O����O���Φc��_@����;#O���%?�U��޴B���`И�~���D�lA�'X�N��'ᔏnv�q��4/�d���ş"e(vgX�27���?� �O��@��KCy�'L	��r�B<�\@(\�t��dJ+V�<qQ��O��4�����O�ʓuH:�@j��ɱ�j�,=ݪ,;pc��Q �v�'T�{����_�������Ӧ�Ŏ��ܤ s�oߒm.�9�4S���
ͨ�6T�V���<U��;`�֝1
Ϯ[�>O��0J�M���K�X��p!f�'\�Dն!g�6MQԟ`���\��:��O�Ĕ�#M�@��$�?|dP��ͅ(��db4�'N�'��$no���O��lzމC�%�4m��Z���(N�(�Њ���M���i����'Q�Ec�$k�4�S��$�:%�@0� �P��Ǻ�� ��_euY�7Ot 	����?)������I��?�����M���'��R�oX	O>>�zgk�r���
f�'���'��^�pz�aZ�b��I������ɚW���eI�1y��ڵK��"�^��ɫBL\�AD�ɻ�M;��i�p�)�'W�h�ƪ��h�n�`#�5_7Jɂ���NL
��5M�T��LݥU?�-���i��Z��?yƬ��H9�5�� ��5y�+Ϗ|�-��O �$�O^e��m�??�r��d���OD���?P���zfˑ�:��C�"Yw�T��ļ0��n�ޟ,��#�M{��c����ygO�!]�d ڷ�̈J^�He#�E�RT�N��6JDŔաQIݚCA����n�O4��Q�E'�u�fR�؀I �jZ�ޮ�a���-��<�1؏}WX8����?y&犵�M�E�Ol��'{�$ [3b�d��U� /�x�7�G�P#8AI��'h��	��ѫ/$kb�'�B�'�A�� >��q�ʜ"�.��}��e��
ݪL�6D�?)��iT�6��)%d��<xM6�%���PŮډ��,X!�R�oj.x*05f��)� .��AD<O>Ԡ���(X�#�DЅ���'���$@�h��a��]x8ʱ	R�[���{��),����PcdF�C���O����O���R�9����G:O��D�=�l4����dJZL��(�O��d�OƬҧ��O��A���7B@n�ꦵ��4!�r�qƵC� Ph�"�]���hg��_�;㧗�����S�e�E�ǵ<HY��$�<	]w�V���LLTX&M����d��8Q�9Q�`Ӥx{�ß����?�@`��&��\����%��$ѳD��Y`��5㐋�~��ӟ����{�*��O�D�O��d�w3n��͊(=d(�1��?�b�s��K�f+2Y�BHFa�y3%H<6�mZ�j���s%F�5~�<�G�_ןX�`kذR�.yi�bƤH� qD�1g�aU��F3�I3��ֵm�:��C���S������K���?����� FlR�����޳t̘�U�2�?���?���-6:a��?�3f�{3�i��ШGM�)Wպ �����b/*ɣ�'�6�������妝�ڴNy����"L^� H���So�#�N�"���(��f�U����9��5bl^`����<AYw��p�Xx��6T��y�IuΖ�G+W��9�ϵ�?�D��V���a���?�'�?���M�'ɬ%z�zx�*� )th˂`��5�6�<i��ib�ي����N}b�'b���U��)&P��4-�&�'�z�3"�[�.�@X�5�͛�y2��*#=$���(��Hb���q,�2pF��DbA=+�Ne��O,0�	����o�9�?y���?Q��_j�%(��d��,��k2�Y��m��u6�+�CE�1>rJ���OB�d�O���W��'뛞w/�@�بX����GjO�bN����a�(o ~y����6�����?�Ȁ%S=^)��gE�g#��|�" +B��g���	�|U�8O��j�<	2�'����i#��Dͺy����S�sf"�#���%6���O�d�O8�C>���kԶ�?���?��ٓE�%�����8�� 2�?!7JKL~r�<	���M�1��`?��V#i��,��a�t�8Ac6ePG����*e����S�_s��y��B�*�b˧1�|��_���/pp:���m��K�1�ҰS���'��!5S�Z�e��D�'���'�X9 �ů��� �ԓP�D1��'#��i��l�(�D�OZ�m�ɟ��'/?ͻ�8y�@AY*%���1���>b.��� K$���Qg�i%0z���Zq*a��&�yBR�7�^���cC�Ӳ3�B��s W� �tu�7�P51��-C-O|�I.(��po��?���?����|���$�DNYz#	�ʜk��M��$�7-��zWƵ<)��Zr�����'#���Ҕ![���� nŲ�����>���i1Z7혶��d��S��Z��O��4���d8`o�l��t/ u@Ib�oVSD����'� ���������?��d]˟�5-T =��� �� H<�|˵�i'�q�rX�������I����'��m�����H�
R<����`���H��Ќ�y�e�������������OV����m|d��"Ο�	�GS/Y˦�x�B�S��� �!�F����_/T`�^w)$l`�(D�<1_w�~����@z��E㎖4h�<rABY08��T�c�w�(���џ|���?���DU�sޡZ$F�͸gFIEW p:��jy��'J�ق�Il����M��`R��vl�|A�n�jbL83���RH��@�F[Q?�0gI�mh��i>a�ҡ��1&j��aK{��;��KV�Π����L;����.�;.xUh%�'�ӵ�<�'�@i���i�J�d�O��$׀B�΁x4@�9��%XsL�^2(���O@�n��!v��?)��?��'aR�V��%��(�\�H��q�eHF���$�yy�'Λ��~bi)�@��'<"伀���}b>a"/wc����M�&Ӫ��6;��!��?A[s��O>驓��\y�bF`� �"�.9��1%�ζ@%��$��\C�S�O��4�:�$�O&ʓ:]�!$�hš���&�������QUj�4��DQ����	))���Q��	!�M[g��^O��F�J&-Jb�j%�H�es���	#?�T+6�64��Z�'�F�׺sw��~F��ɤ6��E:!$�;*.,��S�Ӱ|���$G�����ڦy����?9������]����Ԥ}`�;E&"�9eDH,��}c&nL&^ D��O������pnZHy�v��Dz�.,Y2�6�T�S����:���m�5�Mk�KC?Q��S#]��9���?m��Ν�9u(��G�/� DZvA×^"x{c�ߴ]���ɥ<��ɵ�'hy���<���'8�D���i�p�č�wP���j�|<s �آuT����OF���O��X�t��Ϙ�?i���?�E A�%�z�8�"U� -�X�P�ݥ�?a�{~���<���M�e?!bHѬz�Hd��I�!g��5�ӯ+,�s�s�r���*Dck��1��`�*�T,b��'+�����u*�4���\�uv�+on�hF�'���'��񔢔���O���'�b�R��D�:qcW-"�=�U��*&KR͍�4d7��O�����}�I�71.�Ӽs�(ۀXZ��c͆��pY�'�w>B}�W�ԛ��ϻ5H(x#�Q6|�PY��'��8P��c�M[�.��+ǔh������<N✀m�<0�'�����i0����OJ����NtQfD{�r�arg�����CaLܳ=2<ʓj���Aa��(�?���?������O�͕@�cf�Ш{ �U�_����S���FbӮ�3��O$) d���iN�4�� H���L����
D7J�� �,��l�[v;O���]��?�F��e9�	��?Y��� Q�ubcS����x���*��/�?����?i��?)(O�0yg�#>L�dv���)��C9Tސ���.]�#��D�ئm�	;	��9c�	�MK4�i�B�K���.�N�A�[�;tTA�Ӌ��I�n!�j��=��X�u�'�d����޺S���+���	��c��wd�$z��_:�x��2��9$(Q��A�O����O����e(D���n�s�Y�UD���ݞ.~®���OZ��(!�B�nz>=�	�M��$'<<�n$Z��U4	���SS��$�LE�V"y?���;h��ߴ�ZG#ί��UE�^�?���̡r6���a�^ddɤ͔#�Z!�W��O�I��Obyrg�Ob�@�~����ԟh�ɹ7"d����E ��\Y6��"%{ ��I�Е'���gȃ��R�'^��O�.6m
\z􉄈		^1�/��j�	���$�˦M��4�|���~mӡ�A�?��-K�C(Pef޾a%,}ɔ+��@��Sˇ�Uf[XV���;S���:�*O��-L|Y!pn��+�P��׬D�#\����{�tx�#��Of�4���d�O��U�ǭӑ]��)5J�4t� �2��B|՛��'���q���$�>?^�I8��$�`əd͟�f�!sMU�cA��ܦ]񣢛�q�moO�e���I��������C�Ú��y�f�G/�h���B�^*��� S��?���'~*��i}V�D�O����8P���|���?7\��!�-Jo\��1�J�:����?���?��'81��O�rAd��x��I#�í��TJ�k۞e�H��	��m��ĭ�HZ��2P���	���%,��eQ�ir�kH�܈��čs�B��� =|B�$̆Qtv��'�p��w^�,���n;L(���?Y�P�-%�LcA�+$����`�;�?����?I����G�&�
�Ӡ��O����O:��c&�������oR�A��O��҃���Op�n��M�q�[]?)fN	{r�ɑ@S�?8>���ŧ�ܸɑn���������r�H�r��'0f�ΓJy�Kǋ
w|����Hh���� �B�'%���2Xq�Y�����'h��'N,Ě��^���+�ςR�)'�'�t�S
y����O�\l�Hhp�<?ͻfErY�5��(t�j�Ch3�h�kf��*�b �i�}
H}���jѤܽ9(�%QE&���"�\��5*вD*p�z!F��&mР�����˓j4B�7[s�VA�O���OL�Iʯ'*f$*�aB9x� %��Z�[�4hI���<1V�˒bV�����?���2������'����e.6'Y,EY���9<����>�v�i�h7�C\"�d٧s\l��OO�$ɜ�Ilr�p�W%�z�P^� jD�dYp���i�y2dO�N����}Ѡ�i.O���,W�8đ�F@79.�s���U�D#Ƈa`<�	����������y���u�6�� �'$|��#�8J�2)s�!H�re�'P7��Oz 1���H�O�lZ��M#�#�.=?�D��Z��m EBͼx�"��ۣZ
����<��'�,;���eu��ZZ>����_���5��2]��cj�B�@��G��?����?)���@�����@b�]\�����8am�ؖ�^��?���?b�oe��Q�X��4�?q��V�<��@
?����p/yB�h�o��҄��?;��ƬO��M�'��%`a�:$�Γ����1�C37g�r�S4u�b``P#��.����8��'U2�D�e�6m����	Ο80�&o ��3�c٘M���ib-U̟��Iry�# �Ugh��0��۟�����Mr�/� �:��bZ�%��U}~�B�>���i¬6��#"o�D/H��(�O��(�P�L��Hm;��L))o�٘G螀��0iT�5@	ܨI��J�Iџl�E$�����B�%[6H�a��4=�xd���2a3�I�D_��������i>M�����'� sp(އ9�^<q��Ċe֊y��5;��7M�O��D��Ic�m��I�M�pnS"l%\P����-\�<P�d���8囦��x��ȌW�n�ښ'�`�8i�ú;ӂ[�O,��(3�BE���ǑQ��xJ6�QVG�O�]��n�&��	ϟ���?Q� �Q�t��b�fy�F��(�Q��$(q��˦���|`�	���ӂ�Mϧ�?iE��y��ϟC��D�c�K:�q8A����6M�Ӧ��bE��d�&�V#@��_���CKX>!��͉��*\��!�ɨ(y���d���2Mǝs������ʓbsҎ�'$J��<O��Ʃ_>g�
D+����B��'�jaQ��\n�'��ɲYl`�t�M�(�Gi׭3Y�$ �����n}�h`Ӯ�mړ.u��ɛ�޼j��%�����5�)\��5u��Z1�3F"څk`U>��2K�O���49�9g� *#% gN!rbDm�<�Љ)r�t��ብVF����~���v�=|�I�����4���릹���U���Ӽ{4��>E��Q3-�Fҵ�_�G�Q����"5қ�(A>�^��7Kܛ�0�!�'�T��G����d�� T3wGF���τ���[�H������Lr��ԦU�<�'(ʁY�*@)~�w@�$�$����_~Rj��� ��"�'I��'���`���"T��!����/Ss*���e���J�O>�nZ�M��!@?�1�ުS���g�i�E��*��<�v��FO���� ٓG���K���<Y��	'?	���K2���'c��d�$/�̀�"�^Z�\!�GB�5P�Œ�d
}azB%���
t�'l`;����o~`:�#F�,I�'�6��O��0����ON�l���M�p㊉_Fd!вÐ�dS��
�	��g� �ð�� 2�F�8���<Y� �PEv�$d���P>}���~�J�0�gP~�PH����<]�01c�����Mk�y�Oǈ0����3Qڔ��
H�2 �
�a'dʓ�?1B �;
E�ΟАnӟ���w�����:N�)3Gaͩ����d~b���'f�͹1&�^���Om���̜xy��j�'x.��e�a��Z�!��L��#.J��I pTt�h,OF=��=^��UmZ;�?����?�EW��"���Nm!��N���?y���DϨT�He�g��O����Ol��禅ڴd�9�4�b�j2������-?Q�T�@�ش`��F��~�I�aH�}�g�? ��`D�� Q�8��,J+y�Ńp�J5*8�GɳPz�ܡ�8O��́��?�e� Z��	�m��1���r�49���˲�D)���RG��6���?Q��|2���?�(O:9� X'p�Ah�i�A�5��/��l��ɿ�M�S��0�'� �cћ`�n����f��2D�D�Ka�6�� ���@���m�t�1O�4� )�u� ��4
�̓k�T}b3�L�V{tt���l����	�?��oT��M#��'���'����	5,��ӲyWt��;̹s�g
�7��4�%`��\{ؽ�I������?����|z�n��w��0�a@�M�e���O1����a�8	lZ�@����6Y� �pԞ?	��6&ǎ9��9�bh�� ��Q��ŹL�
h���	���;��'�l�avK�<	P�'�6X�r�i�@���C�N�9@�A3�V�ks	7A6~���OR�d�O|˓d*nac����?����?I��=U9�TR�N��y���y�H��?A�EEy~r$�>A��i��7-�SY�d_*9�H��3��9U���S��c>TK����y2?)f$@�0��@(� 9��'�$�].��F=vL$HQ�ʘ�
m�1���'<R�'z~�:BdXz�OR��'0
�
�ܐ��	�)j�o�,?]"KD�J�6�O��$OԦ���k{^�Ӽ�%E�Q2Bl�D�Q�~���D��]��A��+K��ϋ]*8�J�o��b�Qs�'7$�Е�Ӻ�R͎He�9��$C�=HblثS�V��P&�<���'��@�"�i���$�O^���@ڲ����bq��^E�u��*ߢx���{f���M�?Y���?��'Oܛ�OI�M	 M������>����]N���P����s��[U�O��Ѧ��������rِ��D�$��٘!"׭Fw���0��f��� t9O~�(���<�?fK�0@C剝�?	�F��sFFa�6��+�m���0}��.��?����?����?�/O6�I���6���G����`���"�!3V�Ķn���ߦE�Ɏp�8�n~�ɖ�M#��ie�/��}��ߊMwV�Pu��!1�d�xƃ��.�S�I��y2j�g��Y�;@�$I�E�|���w��Ԙ"ielm�M�y��c���!���,�O����O���Zqu�����EV�(�-ܽr(F���X ��D�O��$��G��nz>��	>�M���/,L}�*C��)���k�1ش�C?l���"�E?��H
 X���Z��|���<j��s���<�RcC�p���E�y�����EӺ=NR��/�OZ ����Yy���Ol�bc`w�N]�I՟��ɣ5��c��5)<r�H�d6����П8�'3
�p*� @��'���O��6m�7�:��$ @�H�v*n	q�5O,�$gy�'q�Fɇ�~�'�7 �ɐ������MY����7l�H <s�<U���P6]�B�͓�u�`��?A$䞗P��I�1�0�-YDH02���?bT`8�K,�б�FP��?���|���?,OJ̸	a�hEj�)L�pH"y�Lߛr�b%l쟬�I��M���N|���?��U�Dl��|p\��2�K�n�p�)d)W�<Vl�ߴZY�I��B_�p��{��@8�?%�P�\�]�r��Q��=Od8�������1��������'!b��7^"�6��ȟt����T�
�R)�O��h�%-��+�g��!D�h��ŗ{��@��'x��'��d(|��I�O��mz������kސX�FlX�ۀd(R��M�b�iU�Iz�'�8T4�p��l��%S��(�l����q� 
)!������'��e ��<Y�� ��D��@1���֦٫��V�� %^[�j$b6�+<L����?1��?1(OK�4��Q��'B�'����H\"���Ĕ�T���d�'Y�`i�'E�,�>�c�iҨ7��)-��d���P�[��Q<Y�m�'gK*���̑�y"`Z�@�&1���.TƊ�{*��|��0OB<��7�D�wDRY$�Tx5I�1+�Tm�I؟p��)UJ"	j���{���iމ�$�Ahm�����"hf<}��%�������ܚ�Ms���?�g�ikRo]��y���y �Tq�a���*v����A�j ��Q��7d��7M�"k���I R���8O> ���u_c.��'�@⢝b��-�;d�ە|#��?B�	��M��'���'���	O*0iQGL�'	8��3$��n�:�2P���EY�W��}���� ���?�1��|Z��[.J� #Ҽy��e�5��p�R����4X�f Z��~���	���Oư�PD@=/��	�)�ѵ�_���F?�y�@�"����I�R����/Ov!���zBr�2� Tn�l�˷�	&lQ !$Ã:_vm����L�Iݟ��IJyR�&N�"4�'��#��6}dZm���ҾT����'��7��O��W��Xz�O@���O��A�IҪ2�(1�W".]ٲP��CӅ9�n�a�M����ؠq5O0	�̐*�u7��	:�tՔO3&��O����.¹;�԰�劷��\�$n�Ph�	͟p���?�dƇI�s�ѐ�ݏ,�^���%�I����F�͟��I̟��ֆʸ�M�)O*Pl�͟����w���\�����T(l�(��d�`�t�I�aN��#E�O��L�z�	�ŗ�J��
�o��*��gɔ�
���&�f�2�" `�rR�N� 0���$f=:P���(1���@�M�b��v̂#1���d\?'�@YA(\Z�􈳰F��2>��4�@uYT鈷Q&��A@U���MRqض*L�����*��4��Go������	���
Gi|`�B��9��H�
݆\�UE8q{� R�>ߔK�E�>z0�� ��}xȅ	0��n��`��v��:G_�
�Da�gN�"�����E�%K�D[�P��`��옒�
�27gW.<?f���8�x� ��ݻv���nZ�h�I���S�\P%@�oɃL[� �&B� ո��N���3W#�O����h� ��.�����Ӯ�0�uqf5"|����ަє'f�%�5x���O��d���'5B8�ŧ��4I�Ea5�Ғ�t���+J�M}��'����$���+��O<�HSCD�4�Jip��Zj��h��4*J^�2��i5��'�"�O����r�͓qj��Q�eK��sT��`Y0��e�i�� ڍ�$5�1O�ca�,�$m1b	X�}�1���ަ�����I2�FxثO&�$3O��G2q�f�ۣj'$e	���-���rSe��M�O>)SCגV�O���'�ڶU�PI�v.ʟ8��X (ҢrNn6-�O���$R}����yr�'b�X��q�? ,q"i�Dc�U��-�Y���a�Q�c�H/�ߟ�����̖'>>Y��.K,8Z�i(�ꗿ��	3�m!��Tt���?M�Q?���L�I��،:��(����:����'�i��Ɵx�I��t�'�l8���>����[L�yEK��Ĳ���zӘ�:6Oj��\���OMB�'�nd���O�Aw���� ��Ӑi:F�g[�4��ߟ�	y�.T����'�?IwG	�Q�T�����8w����4#��&�'�� I�'&�8;���?Y#+M���'���˔r�^��bONV���y�4�?�����X���O��'���	�CB�<h�k��@��HŊ�'������?AW��w�'�V�Q�0@*�%��"-�Xf6-�<��(���'R�'��D,�>A0E"\N�9D�ΚT�D�M�)�����?A͋���'�ܓL|"�L�z ���>G��9�sަ1�T��1�MK���?I��rp\��3$���cw��%��t� GyzXi Gm��M�����'�
�K����'�
-)V��ny��É�N��h/h�����O:�ď��p�'x
���'��A��M��HZ2EC�'�� �.%�a�B�%��2L>����?���i�RDje��7�Z	�LY�/ND��i�B%'��&��ş�CO7񩚧a�x|��郕 ����W6E�'-bU�����4��UyR�ĶRtR�"_�2�ˑ.~�ZWCM�z�����d�O�!d�?���u�̠�a(9W ,�S�e[��Mk�����O|���O�ʓ?\Z�+�1��IK m�s)j��G)
/-��hP��'�:x"��?�b��f?�Syy�ODBBZ P8�G�W;�D��e`�A�~듲?i���?	/O��b��Hh��n��a��nϐ��M�n��ْ�4�?�a�I?����my�O�����P/?4��ׁ'q%Z��Tc�����'��I埠 B��_���'����5�<N���Ā-XO,��E��8���I�bPj�Dl�����b�DxZwaR5����a���K�y
�%+�O~�D�qp&���O.�$�O
�I�<i���8y�N]x0�E1�F����&J����y�曤n�FxJ|�"JߟZ>D�:�	�kv��U��u��B��M����?���*Z����8���1�E�!�`!�n�y��	�T��OX�R��O��?��?��ퟘi� �NBܚbDK�ڴ��d���M���?A��&���1 U�P��8��� (�v)�,��	c &�6�������M�����9��3?���~	B�7K�,���/��@��>�M��Z��-OĹ2���'3���O|޸�ѣ�$Q`�X�� :��g`5�V��1O��D�<9�v���
�dd�Dͱ�c�	`�x�C2*�1��ݍL��$a�Lj3�O�t�'�iF?x�#d$%/������� ݞ��d�O��i0RX��`��A>��ĂG$tZQ�d)�=0���ǚ�?9!�T���ɚN�@��|�-���D:���G��-7�T��禎?R�%�H��Oy2�'"t!�Z>��	~�����k_�,���(�Pڴ�y�CYH?Ѥ��ɟ�Ot��N<	e��2A!�VCs$���K�˦��IԟЖ'P؛T��~.�M����j�F=�� 0� ;�|(ҨG6M|iΓ3�@����?� �<K>ɴ2�B�
��f�8%��	+,Y<Ղ�i��I�>����ڴ�?A���?���+Y�	(]�=���$A���E�%P�% �.��H�I<���	������ѠG"�逿ma�|F��La��m����ܴ6�7M�O���O��}}"�P3�y.L8k�&L�k��h��	��Y1��6M�1s��	vyb闉�O�b�W�f	�mS���$c���1�Ev�6�O(���O�Ӓ�Q[}�)�>�y��'�t2�4<���L���𰶠G"n�P��'d�	'W�$��|"��?��>��5�a.�-b@�36P���P@��i;R�ې2>`�P"I��?i1��<	���1�\7�,�ұ ��,7��Pq��J}� T��y��']��')�'��ɤ�K�`X
9��1���ҵ;�^��������9WW��O^���7O���O���	?w�|j� C(?l!P�䌖��������ןd�Iڟ`�'F���.o>��,^�B��2��
&hUI&�Rr%�ed�|�I�}�\�	�?����%v�(�WG	;L�S��KA,Z�i�-M-�M����?���?�-Ov �7,T`���'[�����9�N�q�l�;N%hq���y���$[�a�]���d�ORAP�;ON�4���	�$]ZT)�д	�
��MS��?�*O����EOn���'l��O�t�BM ���2�
^tb�e�V=�yR�ϑ7BR�'�<0�'�2T����wk��C���5c�h($N��@<R�4�򄂴.JhlZ�������S����l��l�āY�68C�
Y�Ob�T2$��O����J��O��R��$>� �eS�`��\B�bǵLq(�y�o�0��qئ��Iޟ@���?A�O���g0O�lR��¢���hG�=��}q���Ѧ����{�̔'�BA]��O��B�����G���|�l����6b6�O+p�>�Ů}ޘ��'t04�'I�E��M��P�+�0QQŬĚ^����FIȦ��fyB���yʟ8���O���P�B_�AQե�3P��Ԧ2޵l���b��إ���\�x���O���=O����t�1��D�v����@��R��s(q�@�	͟l�I����IDyR�+�����BZ96.@��3F�MTm	�G�>1Y��	˟�Q�	w����؟����q����b$L���9�꜔;+$|�ѯ���'h"�'��O2��pg>���� |q*XӀM���xӆ��r?O������D�����O�xR�_�� ��ju�\J����DJ4^p��`aZ���	���IKy�"��ot��'�?au�T{�� D��*]t�������v�' ��'��{w�'�� ���'��s&�M�hh��M1d�Xis�4�?������"���OB�'�����=;���2^�HA�K��k�5��'�d�t�'��#�O���;62�I�^�'�H0e�T�(
�Xm�Byd�	a6m�O���O��)SC}��F ����@#UF������c/b5p��'��Cʽ�yҒ|R�.��')rh��͹kJ%�8mK��nڃ 蔨"�4�?9���?i�')���#GK~�	�@�fX�6�	0?�h�sΛw����4adR�ϓ�?i+O�����)�O�bd+�uR�17�5G�e22�����I���I3pH�  �OR�26OX�d�"Hd�͞����0�H�<u�� ��M������yZ�?Q�	����ɥ�Hs��`J<�"@��?E����4�?��F*���ӆ�	����fg�,�s�QR�eN�:HdM��&�+G��`1}�L��H�O���Od�D�O,���O�˓z���X!X\z�
�gC��<YQ���i���2*t���ʟ ��s�,����Kb�sՋ��O��,)s�A�}}*#`m-?I��?����?�(Oj!�p���|rc�>~���"P�O��f����7��5E+���O@��T7O��I�O>��صV��d�
ͨ��sRn�쬉'a�-�x5�'�B�'�[�D�I�'����O��K���l"u�����u�z���Z�5���;�|�	/0BZX�	����w���i>7�C	I�z�+�߁&U�5s3�U����'��T�`(s(����'�?�'A�lx����D���Z`�ʐF�\�&� A?�M�0�ɛY���c��7�yw�H�qh��R�*��b���M�,O�DI�K����Я������������M zD���� 8�.�fJD�)�l�IП@�m�џH$��`�/��щklJ��g�L�	0q�U(F9�V�O,X�6��ON���Od��_y2���<��F�`)�h�CÎq��y�]� ����?[�"�|lP��O�o��W�l	� /͙z�:Р�j�L�7-�O����OP�{��zy"l��<I��~�oZ 1�,2E��.}wr�w ��7-1�d�ON!&>��	ß<�	#�%Ґ
� ^��j"�8GD�Jܴ�?)�k�&N�	�e&���O�`d�?�X(^��0���0V:t��tgQ�s���@�<Q��?����$�-Qq��J9��UaLR�C F�"�E_Qy���?��u��<�O�2�'j�@��$�V�ঀZ(�$T�b���y2Q���I�,��Dy�jϾR~�S�#�BW��Y�1�P�ۂ����ɒ�y��'��������?I2��<	&6y�L���왥E�H(T�ۆ c����t��� �'!" �0�?�����E��Y<�K�P��u��&v�\��-w(�DX)k��'7�d��'��kvX�'?}�d�CX�_@:}n�ß���lyR'�Ӫ�����VX1�lD�D���UdN��L�ъ��r��	 C��D�O
�y�M�O��O��;	����J�B���	ܱV�o_y"��&k7�7��x���'`���<1��RdP��PF�*l�N����Ь[�`�I韀��!�x��U�b-&>��p�5 t�w�4���J`�~8yU�[������I�?��-O�Z�'� h�V� &Q}P�s�lГ:��%�� |ӎ���O��OȠ���I�O��CAU9��ISu�k)��w����I���	�p�HA".O"�k�'�(W9�MCVN�������t�Fd*�R�%�������ħ�?���?���=PE%���u
��q)��!��F�'�f���Ϯ<�S�@蟈��:i}������>6}`H�ٙ=�u�siJc}iR��\���I���	sy�L��h�ly�`Ξ<ˮ�'���u��<�%
�������Ty��'�?y��^����-��2��c��%&��r�A�?1+O.���O���<a��X�_t�V&r�(�:á�9\0���*`r�I�<������?��	֟��a�՟���҅pW|�q0i�?$nT�ڄG�����O����On���O���OL�D�O(���T�@8� �iX�BHu��H���IF2��	����x����4=��'��S��?�xU�q�L�2>N�(�4�?y���d^�>�&>E�	�?�S�פd�pq� �r�Œ�=��dZs��<�T�4?�T����'�4�]Fe	8���3;�܊a�6�&6��O~�DE	^7v��O����OL�)�<)���ƨ��N
�h$�L��*K�3�xi���yb�aRL�DxJ|z6ū-�	��zin �$e�ȤŃ����̟��I�?��Пب�p>�yUoK�t8�)smΡC��1WϏ��?	�I/M(#<�|��P� �aG�R8�mJ6_@,�s�i���'b��%�h�m�P�͟dZÍ�9�xJ炈�F�<��&�͍l�F(I�}ZXt;�yR�'8���EQ\�@.�E�@i# �_����'2���Y��z�p>M�I�0+b��r�cC�22���A�@�k���if��x�>)(d��?��?!/O�qj��XM��co�j�h�7h���~(�'W�	���?ya�^q�t�'c�,G6��y�Ey$$���P�:6Kȉ~1O����O����<!#f�U$���>'�!�iY+2z¥pwdB&J��
�?)�4���?�	���p$�>�BԘd����c�>[N	�Ff�A}�'�'R�I�m&lkJ|
]8 rc�f<���7#����i ҍ��~����?	�gh ��>��"" 1tm��_)�V�`��[æ�����'���A�c1�	�O��)�7�i2��Z�d�rH�q�7�j�b@�O��'�gS��Oj��{�? �!QA�&��;D"g�E�&_�d���qd$�������Ɵ���fyB�ū	l5��!�T=�0ې���KLعj��'�D�>cV��A����+T�pc૘�'�f�S7*&�M��#Y9�F�'���'	����<1!nF柠AE�ޙ1��H��'6*!��^-�?9m$�O�D�).�:&��a��EQ�6Es�n�����O~����;{@͕'ry����?���O¦���2�J��τ�\�2e�p-+�	�nb��Iퟘ��.sb@�E,��q�`�U�5ZD��4�?���E��65X"��Of�yd�?טq���!U.--!B��� �=b�F�x��=�� ;�g"��@P�Z	t*�:��
�$7U��'�0����vc��;c�-���ڌ�d):���[G�ݿ6M����^�D�����0h	�,{F�I�S���	Co͛;4��#�̹q�����+��>�����&DQ(L�ĮD�g�*XH�iLv=��)9g2-�.��4��b���XA22��	̺��`�Э �r]a��ٚ?����+Ő5|�9���
)ۀ�Ca��s� 9X�Ne?L[�L:���8�+ƲR���'��r��8�̹0��NL}���R@I���8	�=(��˶���zc	H�'�>Pð>d�	!d�'�S���	���;��q�Cɂk�<�� �Ɵ��	R��R��@��(��9= Dj�(��_]H�ϓ��?I�^=q1��J�r�p ���x}�G2�S��_��������!���}��(j�a1g��ߵhڌ�2O����|�e�A�?���?�Q��L�l@��@�K	ft�K�4�@Qa��G9/z(���l���b����@��'��#'(�$r�B�<.,�0 ��i�C)M*SK���"�O?�� |�ލ��P5�da�LF-�����Od��,?%?]%��!��ve:�)��?9-j����3D�|�o�Hjt�����H���7�$��<�Ts��z�'Ldlxu��a�|��	�@ ����'B�@�����?!���?ɨO��՟l:�F�I~��i�+�a���Q������ˁky~�j��p<y��ƚbd�a�(�$���ү^p?9�E@�r���x�JF�I��x� �
*���V��f�uRQ�O(�~R�F�?����hO�ʓQ�b91MD,5���ض�F�-N���I �yiܭOG�e�ge�DX���Ї,n8dX���O��<�a`�kb�[�U2�1�cݩt�vA9�@)���Od�d�>!��$�"�'����ϔ$.��ם���8Q��.^�z5jp%A7s����	?��J
�q(�!�ʈbb���nNP�\�G$�<,{r<��I8����Ojq��] 0g�D����:��p-զ��IYy�'��O�ӣN"�D��d^���9��Iާ
"XF}b�#�X��3%�AIPL��H��Oz��͓GD�Q�i��O��IM�B�r)�RV#A��"�+�:�B�I3
x\�CFY�D��iI�IT���B�I!.�C0�������fe�K�B�	/}��T�( a��@Μ"5ˌB�	�a�ƅ`��',.4���+�-L�PB�IN��GA�V���c��0[�C�I�7 ��H�%C�!�|p��4��B��.c�C������	�*C�\]rC䉆kU~ 8�C�[��|ʥ#�I$C�ɋtgx(��C�P��T�@�T�B�	6}��H��l�b=�̫wEE�`��B�
(���! %f��x�4��hƌB�\N�x��O�t^��a�^ XvB�I�	J��ЬsC|����:��ȓ��`�6JM�4\�51A�L��줆ȓ8m�@k�c�hZ����H��1��u����OE�7�ɑ�4�����u��ٰ�Y�HiZ���ꬆȓz�x%��H�^��� ��[�Д��fp�;7kѱ5{̐���M�;���ȓ~�(A[��9��{�$�)����5���SDC�$>�ˡ�P	�a�ȓb�nM�q�Z�F��Y���{^�����A���لW�jM�t%�<`#�H�ȓpb�j���n�h �3�9X�8I��+��zf"Ye
4���6�4�ȓ?҈�"�ɔ�Pl"��ױ\7(�ȓ�� �##�!�D	zaC�,�:��ȓU�݃�K\4V���)ţH�} ���S�? n�y����+Rv<�6&��N�h���"O�\�)a�D�b%^ɮ�a�"OV�"�-/���Sf�,`��ٙ�"OZ���!�6�V���#D	p��w"OD�@l�9g���[�K��2��ɣ"O2���#��13Pz��ͮ{���Yq*O`�FȚd���:�)T<r!$qҘ'���	&��G�R�c�B�>E��C�>]E�������,pyց�,�y2,�nB X .E�@60��j� ;���u!@2��PS���O��RD,F{s�1/ʆ1B~�y��'7Ĝf� fq�lS$+&�d8&�؂Ȩ���4A*,��Dϟ~8�C O\�&�XIQP႐��ȹS�} ���U$)��'Gf��$�0o^,��ᕗ��\�ȓ"[~���n\|h8�� ��=�}͓��U�G���8�QS�"~�t���#S�A�����6�����Q�<���R�	���ʦhҒy����׳_��I4A���P�%k���g�'�d��R��c�Ը��Ьhm���2U�쒤�E40~�y��/a���@eJ0DcČ���S�a��-eF�i6��o���q��G?ʈOD��%�	%�6]�a��U��9#��M:TC� ����q��mO"C�	�G���+��).pl]Ӥ
@a��I�FB���7I��0�O?�-	�2@�H��D���AХ9D��)�bƔ_ˬ�$�Zo�"՝��$�"5� �: �*��3�oj��b.O��v$�
�0i�P8���6J Y�N�<<n�m¥@�"y�2�Ԍ�)��c�$ذ?�s	H�_�h����J�s�:%)!�t�'|>!�rK�P�L|��N:��9S�du��˜Y�<sb��$8%!�ͅ"r�k�����$c��n��$ֿr(��aLL09��է��V�+���R�21��"-����
O��	@�W`Ҭ�w�R9{3�����M��'_8���)Es��Yu	!�C�]2C@Іt�8-�J�a�D��	E�Ѣ4�"!� Ϧd��ܲԌ׸>m!�Ē�P��S�C����gl�<E���`�3�9�)���y J�Ң�B��.5��	&H�fC�I��F��'���Os�Y�/�;a㞌��2�axr@R!4���!@�8���((��?A�@S#0�:"q�:�����*�¥�q�R"�x���yY�}C�H��h��sJ[	��O�E�v m"�c>a�UM��A��- =ږtz��0D���Tʎ�t̨�S/B�Y���<����H�}pO>E�4��5/�ı�%�&J�D��#��yb��/��|���YL)|s�����H!\3���0<��R
�ܩz�!�L`f8�	�y����QS|KBMCw�ׅd��q��8�Ձ7$�v<A��C�n.���1��HX�l� ��P�'5��@v��:@1��(qӾAZ�!��3���k�"OT�P�ֱ/(����*j��s��p�5�+P�tc�"|"��N� �@� uNJ�8M|�BH�L�<�W(�d.�P�5ክo9~yѕ��I�<�����0��#�&�&;�@��l�<A�Ua��Mbb.&'Dz@P�.�jy����$��0��A,��1/~�t��&�9�0���(^�|C�I�:ώ0�T�Y5/)��p��e���$�(�ᕻ-�l='?�hq��-i�`-1&��i���U�5�OJI1V��?�*!���`�D�)w��3�`����R�^L�(
@�`R����;.ja#(�4���)!_�$ ZQ�$S��H�AW`�<1� 0��u�eY��M[&#����
�(�jԨ k����)ʧbT(�,�=QU���1X���]�ȓ}bt`)`DV�-�B�{�a�v`�����>�w� F��4KI~�=�2&7<���a�� fT����CF�<�A�)E`]��Ɨ�n��1EBP�<���'���/�q�Ht�$V�*��3	�'Z�,�"��x�xŪS'��$������� F ��mE;a>���hג
0���D "���OS�X��ާlP�C	�8kfN)"�'�UH��C%U�ܽ3���_0 U &�P���'��>�ɓ\��a#�L�cz}!D��DC�	�|�0��*H�GJ��⥠P)����-��������(��dѿAtFE����1K�{�gU6H���/R��S1!����Ɇ.ܩo'�B�I������A�4y$��⑪��LT��Q��H>�	��S ]�`H�֩�!1�m[C)D� �G�8;�(!t�N6V�`E�WD2x���HG��'O�9j�`9df@	��6`i��'���Re�a�8YM�U80��9=f牛��0?�F�@ Yה���~�4xe@�$��M�r�S�O��u�e�:WY���tK�t��Q��"O��D�'������cY����V�D�vn�l����k̓:֎���o�-J����"�?�O�����~�<���>Is�e/#���9�dĢ�!�$� @��t�ć��W�>�� �]32�ў�˶�e�O�dx���$�1�TNU
�@��'�z5��C�^�4J�� |7�Ia��K6������ӟT?���bFE�p��X�B���C�	�9�$l��K�9vu
UD�a��C�I�h�� $$��"�l���Ǝ�A��C�I�Pl��%d�K^ �x��ΏV�C�	3��a�ႋ&H*���G�g��C��H�!���L�ثe�?�NC�ɍkn�,��#Bt��R�&O�}�vC�IR9��ڧ�K�7���ڦ�8��C䉜'*�� w+�^��u�@��){*C�"v����E�͎Q�n�ɓ��30C�Id���T�U�6G@�;�!���	G؟P��cH�^�L���)�>5~:��`?|O�QO<ٓ���jI�er&
�S����{�<�djW+1Fb�`dh��!���ѧUcܓ8���עA�ȟ�@2c�� N�*���^�b��"O$qBTM�w�(UمeV 0[<��EAUT�sK<!�2�gyҢZ�^x�����. �Pn� ��x�N2Q�\q��,X�'�e�'���%q�'8O��z�[����d�X,��rcնS܍C���#]y�yrkŖ�܌A���y6�1ӿ钠xHK��z ,�4�����'����
��+��l��X[���+N<�)�X6���S�"QN �����c>QpT�ׂ&J8͑b�T�<�
O;D���jP�tG�XTi؞-&N��A�J�. tKs,Ѯ����[$�c?�:�R���&	�=d6�DB�1`�u0Vk8�`� ^�-߆({��??Ӛ�:�a�Z�����e��GI ��7�Ȉg�Fͣ�.�5�$���h8�4)������I�N����׬دV�9�G�	�H��1L�&��C!�9>zx��0�Աk�:��č�:a0�ۢ%0ڄ����Z�D�X�	1!��N	2�sT/&>۴��S�S�K�t���\&4����I�_��C��&?m�yCG	��d������l��.A�w�$���ZV}���Ëo�"���h�*c�R�MAǨk��"�l(<�@�.�8\6��>���ʕ��]m��ӕ!sX��7�	�h��NQKQ�|�W��'m�N� H�'M���f�,,O��:�Q�^Ϛ�C��H�Ot*�j�@HP�<;aG�&^
��̚�F��@� �?�O�madq�m���l	�Ȉp�x�˵_X5��ړm̀�&+���~J?�`��9	�"����Y�R�(���e'D���U+U�c'�,z�/<L���&�5R�8r
ڂ7���05O0�?�D��4r�L.�nP(3�\]5����04��s�P�6��)�� h�c���(�>tE�y ��1��]��j!�_	ԁ�ר��^\%s���m���)o.��y���`6�H��&m`�@'ɍ&4R�:�.ӘGGfqi�X��������KF@T�3�A��q���>�I!Iy�D�S��-��\0�B�A����|���9k����	��ιid"O̘{���u^da��(H�4I�Ĝ��LQXs�UQJ���DӐΑ>�S�? �@��ȠLltcbH�*F�Vy�4"O�q����p�P�/ݜ@�j�)u�'J�|��8qp��`�V��p<��Mꪽ!E�N`�UyׂT~��g����$X�la�a�v���.��80�߰S�!�ǏS��p�ᅖ# t���Gɖ�m�l���7�'p�	�E_�j}��#�u��C�Tr��L4X��&"R2����hO?���ߪmWEIAƛ+/9�YPE5D��w�K5>�ƭP���'K�A��9D�D�p�/C�杙�d��?��dl6D�8#���f�Ā!ې�3�N2D�48s�D�nlQq��4z��!0D� ��ӚIڤ8D���D̄��@)!D�t{��ם�b$i�AW�J�{6�=D��x�c��f�B���ӌC!%s�8D�@��/�#T����cS,q�qGK6D��7*X+l��Xa�K�R5���ta2D��!Q�������A'�:~�L%1T=D����-
�N��<�b�N�
Be�W�7D��ʧ��%N��C�3Kf �A*)D�H0�ɪcLqZwX�H��c�4D�ؒ�>#JZYB�#�������?D�`����+|��F�_����3@<D��p�@�rM������5�jH�<D���a��o"�E�@h��6/L���<D� ���ԼT��j���,�'n8D�hJ1K�q��UP� �zk�t���7D�X���2/@P�bF!ߓ"o��Є()D�4��*p�������fR6��%(D��V)��c�����3U�h���#1D��!@+͖x(Y�w��>�L��3D�$�$m�@��4!T+�/^��]�A0D��G.�Q��8�Έ��4��A�1D�pIĀ�10m����e�9*X$( ��0D�����C+��"ဈK>��*P�;D��y&H��W�����J����]�F	7D�l�����v���#Ą�%����:D�����P�#�#Xo�x̃��7D�p@T�: ؈��7����"D���M��⢉�IP^xXӧ?D�X[5+G�?k��"���`�py��N>D���Δz��p���bQ"d.D����$ϵ�Dq�!߈v{*eiEa2D�`
2��Z�=PPI1D����1G��æ��>R�|�3D� �k�UK���هc0�;�D0D�X�#�<z	�ѳ���T$D��h¨�cn�Y��yj�Y���!D�)5�۲���BȎ�SѪix��<D�0��o�l����&�L�*0�]P��<D���F��Z�rM��ġMV�����;D�8�J�X��#D`��;��|+d"$D�d�QfT������J�ļrFL#D��z!�:Ph�ʑQ��䚒<D�D��m�J�x���kr.�
�%$D�\���Ƒ% �b�E�(
A�����<D��h���T���ѷ'�O�T��?D�8;@o�0eO�@y㈺uj4#>D�L�"��/�p����6P�P�j�M;D��Rw)>v�]���auv�kq�5D�0�ˌ	AZ�E@�S��:<q!4D�DȱMA�|аH�T'�Z�r�1� D��{D!O�TvΝ#"�˸T)3e�*D�Ȼu��L�Z���?Ge�șR 'D�� �zQ�B�K���p�(��B`T�0�"Od҂��\v�Ç��V��H0"On`� �7$qX���@mT0�"O✲�j�wXt��kIRL���S"O�)*��Q�#1Vmń�.O.y"O�8�QlK�fi|,�NL�X8�� "Oh�b�	�QY��s�GT�YH��x'"O��8^��`�����EJ(J�"Ob��tn��h��i�
��	b"ODɀ��<7:QarGN�1�"4�"O�ɐ�k�;�^T�E^[}��0"O�B�I[eD�Xd�^]�4�P"O����
�H���d�@�#$���"OZ=r5�1p��ԃ���(�"O��[��aX�T���*r�y�"O����fG�^�h�@���^qZa��"O���%��4QV�/��<���U$I�!�$��%�l��A�A2j�̴7Ň	5�!�$@05n
�V�t������!�E�*�j�*&ȑ�SF���S�4�!�Okd��R��&2JNq���Ɍs�!�֊�Pt+ͩCA���-�C{!���3T�|a&��n^|	�e�� X!��Q�C�,�2̘�KQ�!Rfů_!򄓻2�x�g��K�h�%��4ia||"�7zq��U���A�l�'�y�?.�����.�^�����y"�U�9�`�s��J6mx�i�F��yR�L�T�	�@��- 4�c��y�DU�X4B-��B�*�8qcP��yR0xe.�iD��9�"J#���y�]�P��	B�5<�E����y��B�h�B�9@�JuЁb�?�p>!M<i�-��6PիP�Y��a�h@�<�e_�b�%����!}e��r��Vp�<��J�X����˝H�$�`"�V�<�\#0�"d�A�$iv*ʠ�ST�<� �gl�t��H��xL�<�co�:tW)bF�(G?ɢ��H�<�U�[��%1v@Z'm��90���E�<&��48�TA22%�t�aB��j�<ɒ)�.���o��
�P
)e�<i�I̬J�L�ۧ�\	V��u٥e�c�<�Õ� �2�!�����ҁO#z�B�ɍ'�#�	�:�0�)R�˚zejB��c}&��Ѐ(�P�	�K�1"�2B�Ɇ7$�3KZ�7T
Ӏ V��B��	v"��"����#-�B�I���swD-!�u����u�B䉃ݼ�#",	.D��	���/D��B�I�'�L����\���B��
�^G�B䉋p�Jt����T�,�1�̥O�vB�%'� �-�C.l`(fj�-�B�� P+�q�UL�F�48i�'0G�B�IS�4�!hْ-���fغn0�B�I�z0��Ƌy"�c��$anB�	3[�¸Y���
� �`qC^._�LB��#C��X���6G��H�w�^fR�B��+9��rȝ%kv
(���}-bB�I�~&] cm��:}��@î�}>B�ɷ�~)�faĳm�~��hW�mjTB䉉xP�&J�r��TA�QO<B�I�=䄽1%ĳ���ʜ9V���DΪɔ�a��,±w�!�� �����_-6�iC�Y���"Op1������8!�F#5���`"OR��$
�4���h����Q�"OA�E�-
�p��ϊS����'X�O|�V��	�e��-�*\����"OTIW喿��-��S���"Ot2U.��|� `A-� �.�07"O:\��o�jMr}��3<��sp"O�(��	^���ҧ�}��"O�@:�}��S%Eo+r=t"Oz8v݋.�ʄ�T���W�٢b"O�|x��$�LP"ʇa����p��d���I��ED"5+!�I�yg���NI
!�dъ}8Hd��cѵwF��p��|�!��M���d21��%gˎ����'�!��S�T�9%gؤ���"h�!�!���[��y�b^�W��u�2��6�!���j�
�%��
F����"�!�ך$�aq�ē?�H���e� X�!�d� 0rxA�b� -�����!��#?w<bd�J9|K������X!���P�^�1�M'O1�H����<�!�Mr����8f#��҂"A�!�{Z���FD�D �0��;|�!�䇤+�xH9��$?�F%*�Ip7!� /h�:4zF�\�+a|)f�E!�Y�e�p���P� B�U00(�5�!�$G.�@�X!D�	xȅq5A�>a�!�d�1Bl�m���Cuf)�1&�-L�!�$[���� k
)�� ����!�#tv���#>�!���6!���I�\9��ٱ	����O$!�Ѣk �w
N�\ﾭ�A� !�	�apr�� &)'�0�S�!�$Ϩ=:hФ	'~$d�s��#,�!�$֋I	�UQ!��(�y��.5�!�+E�p4Y5G���`n�$L�!򤘮0�fh�vǐ�!��B��f�!�D��%A
��늅7c5� -o�!�ĝ�:L�p���sVl��0��Fu!�B�L��������0>��ҷl^Yl!�-|y�S�A�`=�q���e\!�Ò(d 9��5�9�P�5zT!�^;O�2l[7M�����,��#A!�$Z)i�&���E'n*eJ��p&!�$Y�=��q��3=����kߋs�!�D^�B�3!��#��!��`[8V!�SdZ8hg���)hF��$
wF!��׉2+�1�d�$jrN���D�$4!���xxR=z�Mў)L�W��35!�[�	�D�2 Q�I𒍨0J�6y!�d�3��`A��`q��yW��0!�[���������j3�B1�!�$=��9a�V\�v���E�(9�!��iy�����7c�H�"/b6!�[�J��Z�%�\��� �D:D~!��}(|L)!�	:[�����ޣ5T!�$�.D-�	RcY�xTzl���.�!��C���x��_"'#4�ҥ#�9�!�5Ռ�Z" �!x��{��P� �!�B�e2���b�(\C�[�,G�Q�!�A�k�B$��/iKZY�3��V�!��R8�aIp)�x"���/;�!�D�N�h�"@�A� �LjS,*\!�� -��B�� �r5�U^��}T"O8�3r��;}BГ�+ҡD�8�"O�%�*�f@��$�'��� �"O��%�QI��PB���5��< �"OZL��,ȴ&~�8c��1:��y�"O,}�c� �r	�����X�"OV]h�.H,�:�1�d��VT �p"O`˥핞t\̨t��%�
�i�"O�'!X8�0�#"��%xR<�t"OT@����<�}�6��<{<�"O@�(��?}Y�-��D�k[&�hE"O"����P"-q�c�NX�x0�"O�Y�4:�iYFBG1kK�]"O�Kդ��"!�b]�J��X�"OԜP�!�JI���Ӝ$h�IyW"O��id��j��H�7OM�QT��'"O��;0M�T�XQ�.J�}Q1�"O1	U�*<2d�� �3_;�ř�"O��0s���W�d((�Ò9#� �B"O,�����*:t�'��%jc���"OƐ�r�/V\r��g�qJ���"O4�0���#Ez����o����D"O4�y���$���.�,X��bT"O���a��+xR�2�|~�E�G"O���2�kN2LY�$|���"O !Z'ϲ!�%�fO�0b���"O@��.VNH�$.��hy��Kt"O���A��z\x��S�^�Q�&�A1"O�!��e���bmʷD����r"O,���7���C�IC
]�6��"OUqs+İDp � H�6�lD��"O^)�*��t^M�hL�M��@Je"O�Г�-[Q����g�0��7"O,m��K[.R������Z��� c"O�#�Y�0,I
@��<8��0"O���aճ>��8�S��;Ql(�7"O���F
rK4YssN��p�}kq"O�ܒ�&4!Wt���'�}��ecV"O~u � U7S�Ix�fZ	:&��$"O����.z \�Fíq%x�af"O��y�sY>������O�\���"O(�rW��7J(2��mD�b����"O�k���'�H"��'��,�D"O~	�#$�Dl� �`��#"O��a��)B���B��5xHj)Җ"OT�: ��qj�Ꙗ@	c�"O��@4�]7IE�lz�Iɝk;P�"OH��3͇+8r
$s�H_=0�<�v"O��!�F+g�xz�hG�_v���"O�-�6��y�f`��AQ���"O���-D'Z�� ����*�VAʀ"O.I٣&>�<�%��.,�E#"Ox؆��*+p���!*��Dr�"O�����I���|����x�a�"O��Rp�8NN�P���j���җ"O�,z[��-��$�q�yj��	�y�Z_�n���Y7L~�aCu���yb�� |E.��� =����]�y҅F4`��� (^�0�~DQ���y����jJp}�wF^4'�8���\�yBGN2��0;�
����A�`��7�y�(wx�������"U�j��y"��@���Sb
 s�tB�A���y�7h����7����I�<�y
� r�34,R�(���\�j�E"O*DIf��Fnd8&l�	~�q�#"O�5p5�_C��8b�֙Q��I2"O���qB�R� H(��J�P�4XrB"O�m�%G\>z2��E��)�!K�"OlX��f��Nlر NQ;p�6"O��;�� ;N"���� ����"O����p�V �ƭY�u�颀"O��{R��:KhJ�3R� #2Ţ�0�"O�C�0~f�1���;��!��"O��p)_d����"�,�"O�`��.��Hμ�h�m�;�Ƽ�"O���	�%WY�'��5)���"O��S0�]N��!Y���|t�[b"Oz���'�vh ���_Z4 �"O�	�O�љ��^X����"O4�Pb���W>p�$eŻ<��۠"O�����Wϔ��
oް��f"Of����D�[Д��t�9C�nY""O��#����\�2H��%x�"O��0��K��y��-J�D�Z��R"O�}��cɕFx! �L6f�<��"O��	�ى\9�7Kק!�|��"Op]1R��#��x8b�Էy���e"OH�"�l[,Tj�Z��S�>y�u"O^a����#A�5BDj�@t��
W"O��BG�I�4y�p�	5"Ob�#��	���Y'�Z�=`��Xd"O�i�RdǚX9d݈�� )J�\�"Of@)wb<7�T��Z*N1 ��7"OҨ�S�#+���4BJ<@.VT
�"O^d:a�^��<�8�a��!��us�"O|�JF��Y�4��g�~5��"Od��!JV�$` !Ȓw�<��4"O�u;g-��@��E��-�3���i�"Ol�V_�()�^	*w*��2"O@���m\zX�$�J%��%��"O����'_P�}s4HƪTr�"OhՑ'��vg�l&\8'��,��"O��`��nxj��f	xR:�"O�A� ��o�"IF+DP,�"O���S ��ya�D���^�6�*�"O�ЈVkG�)��Rf�(���w"O&�A%��LꐩF�:�nD¥"O.M���ޥv��xQ��͂o�MCf"O��ˡ��M#�)���N�(۔!��"O��)��G$�s"\�
�0Y�"O��cͫu! a2$Ӆw����"O�l3�'Q9xɑ��L�p�(��"Oj���n�6��\�$,A�U<�"Ox L�*~�&p��
� 77(@*�"OT;Ǌ�b4��u(#yv0j�"OX���>q�����
x��:q"O��[đ�nϨ���S�*,�P"O�kfQ=6=Bis�n�hE@5�"O�h��W.L��\<1.!(U"O�Ѵ-�	d(�������3"O ��lR�drvt
��n�2 ;r"OL���F�~N��0�Z��V0��"O�Eb�W�/�d⅃�;�>�
�"O�BQ�4H� @u�A�<@D)A"O��C��>*RA�"�4��S6"O�bce��.4��3�`78�""O��ضۻ�so~��q	eq��S�? ���ueD�6L0R!�_eT�f"O���p�ص�"P�V�M�J扣"O�PA��^�A �YS���;�Z�a�"OQB�4��Q��D;O8�`T"Oj�0N�= 	��)���E�["O\�16�E�Y�5��\#;?(�"O������p9FMO�a�F���"O*apć��?o�,��,K�W�Rh8!"O����De���*���(�z`(&"O �
VaI�u��ق���11s��R"O�)��"z�c7�jn���"O�< %����*�!G,�S�b��"Oe�1w��}yG`Ǝm��HA�"O��jUJL�uA���Ք-���"�"Od �V��6F�82�B���b�"O�� ��Z~���S0	�HBs"Ot����!nK�1UL��w���y��-��S�[x��̓��y�'Zm��CF��~�Pxw�$�y���gՃ�$9x�v�qvA���y*�H(�Y��c@�~�J����$�yr�ߔx���Ɗy�Z]�Wezs!��3y�����`�l=�W�U_W!���<�I����Ski���>�!�D�*\^���@IW+O��Ғ�˗Y6!�d��,^�+t�R�7[�՘�M3)!�D����N 8��B���<m*!��uե�aH�$#�����;T8P�ȓG�f㱠V�xfԘB��w"�Ň�I����d��i4���=hS��ȓ>}nȋ�Aѳn����H� �4�ȓhFD��n�oj��!��<4��Ȇȓ��	s����ߎ�]�R�)�"O�t�d�@5r�T��C�'�B��0"O`�+�m�"Vv9�4F0�D�d"O	y'l�kl.�rLR�3��,�"O�\�tI����B��ϭS%֐�"O6��t�y2�BL�� Е"O����59�|�
��Kpb���'�|$R�E��Ltj��.��t�	�'�@U9 ӌ��Xس%+�\ 	�'�r5�w'�P�M�+OƆ0��'ߌ�B0�
�J]�ͫE�$?�"�r�'=`��(I�W�h���^�4��[	�'#�	�˔�F.(���&)�ZP��'xȱR�K9��:7��&���
�'3��y��HLvYq&�"0Ƥp�''@,s��ڝP��5�%�� �T,��'�h���_�] �������bX��'�D���4�.�S�^8o%I����O�S�g�5dk+1"or0k���)!�$��9�@����pO�݃�/�5!��^�p
��k&��8(?\���c�!����;H6D3�L��LҌi0�&J�!���
"b�P)o
�;���Z$�˰#�!�K�<�l����C5h��䰀� �!�D�'|�u �	����奘;��'��O?��7Ě#xH��
%͋c�ID+Dxy��'ua|��V7x&�i�%
F#7�"��a*Վ�yB#F-�J�B��«FV�	z�$�
�y�������@hNj��ql���y�b����(��@	�+�n�cI[ �y�B�V]P��ͷ)����#���yG��t�^�A�d�j5��c�ǁ�����O��`D�� \���@�&�f�5��6-�R�+VY�|��ʟ��ɋJt��Ɖ�y~$9���>�DC�#<�C+��1DĨ�� ='�
C�	?(L �U�ݵ6*>��K0NU�B�	B�й�L��v\z�g�y&�B�IRM��b%$G�V�.�Xf	��B�I�#�t�!gI#�NY0w-��e����O�����N��.m�C��C�d�*���04�R�'ߐ�f�̨;]l��A>	A�a8�'�n\"@�A Q]�躤�����
�',j�xa/�2H�� ���_(v���X�')$){�gߏC��b2M�?\�a��'�vm u@7PP�R�'��W>H[�'��eZ` ��O���c��)���O�1��0bt�p�iU;0�,��"OH-k1����v掰O�� `�'���A�F5++�<k�+�B��!*MT��g�@J�]�f�K@'Hڴz�.D��ǈ��'��� @`��1z��e�!D� 01ϒe��hc�C?69R�(7� D��;!�:Z�X�VO�kl8uI6� D���e ����HB$��m�2��e D����|�&:�E8��	�?D��R`,�Z�I���A57y�;�<�O�ʓR��Ɂb��{��0!��M4+�*���'=kri���ɕi�#�NT��'v)��G!bs�z�����y2�na�MB�����Р��y��CY�vA��|�D�3m�7�yR�ļ;b�؄j�	p��AB���y"��#D
�%�΍	�(�aT��?�'/��4�X��q	KDV8�
�'�����`��*��0X9V�R��	�'�ԘGd�E@$�ЈO��
�'|���F��LGf�@�NL̎,j	�'1@��j�1r��
HuX��'�$�zt�ܷ���L ;~��'r�  `!K�D>q!����9!�t���hO?I�p�	#*�DL�ǌ-r�2̨$�Fg�<i��98�m��(@����A�_�<�
�x%8���,m�@d�q�<A��� �T:��';3T�ڒx�<qvŋ�8������p��@�I�	g���O��a
5�0��s��)4����'L@�᱇Q%
�f]��0|�"lc���'o�>�Ɉ3�aZ�b�	il����?1C�I	sn�!x�f��[98yS���$C�	�<��Y�倱u<�X �,��R��B�ɢ ���ʒgNf�� � �ڍˤ��$!|��̚��P[e�1B��D��ȓx����&�K.��R��ڙE *8�ȓO��T@c�Ir	.y��n��#
(p�?Q���0|�k�h����/� b�f�IӏBr�<9�E�E�`8+�"Y����2��g�<�T�I�d�01R�i�1[���4 LJ�<�f�6�Hp�vo�s[0x�Ej�Gx���'�JI&�{�ج�Fn�	�p�{�'���b�A�G�L�yW��D��K�'��[�W;J<l�3g�JzH2��M>����?�ϓs�jD�k��T���:��V:#4�ȓ{ ]�%�k�R��"��2�X���EP\|�S���?�(�򱃊�|Ä���}y�2Ox���R:8s��*R/�4:���Y�"OXٻ*9bQ6T@�J�AMڐ�"O� ��D����"����\H~9AV"O�!�A�'q-�B��M=a]@|+ �d-�S��D�(hČ�v(&ycΠ�.S�N!�$U,z�XJP��'	������H0w�!�$��e�qN��@�"��s�|}�yBZ��'&H����o�P��N��*��|�
�'�H��c��b�ԓ�nO�w��m�
�'��C�*\y�<���ι`�Lj	�'w���fL1y�je��*��`�@���d%�6\zueH(hт�%$āa����"O&�P�(�`���:@U�p�e"O�I����X-��s1$k�Qi��y�mZ�p����[#e.� fY��yAջ����S@�I�r�9�����yB�06�8�2('.v<;C��.�y�֫$�$����� *u �(d#B��y�AE�4�n�0�'��G�śSg��yR�����+���>0��dU)�y�����J���	3�1�d��y�ױ�&y"��G�	 �QQi�3�ybie�J`��' l9`Vn<����Z�"�IUΟ�:u4�"-�@;.u��	F�'�p8af�"���O�!�l�:�'W�YaM�ix�����1Qx4x(�'�.��g��h9�x� �XŖ��'�@�V`�!I:`�[��\�D�x;	�'D�q*�;~V��#�,��&I�'
���-A�,g&�[U���7[$@�'��L�w��YL �3iH7�������<�?��%� 
 TD� ��j0E׾]������E�ȄL�@��gףq_4	��ZJP��b��N�H����t��H�ȓ��􁣇б.؆L�Be��M����x�,L*�*�}��<a��ѧ;�ȅ�ȓ|"P�)ñ6*�`$�ˣ2�H��П��	�'�Ļ�dh���Wh�b���O�d�O��=�'{7@M�7D^ 	Hg�ʨo����Ɠq~"���Ԣ}Z��!,��?hBt��'�"�Q����L�*�.�">���'�*A�
J�<�H�m.E'� �'O���U���$�+5剆5���)�'�]{��0X����H��)L��1�'j��pŕIʼ�ұkŗ"}��*O(���O��=a�O�Xu�J�V��|ز!
)?7F9 �"Oj���f�����'ݻw,���"O�5�B�X� �cF͋\wB4�"Ox� �/Q�9��9����w�ó"OV4�bE�=.j�!Ԏ�,:����"OF�;�f^%�h��xJԐӣ"O�9/V:<�Q�=�4�B�����?!��0<A�J^+b�1ڵ������a�b�<q6�]#2X<� ���sâ�J�@]�<����NOx`ff
��*l���V�<��L�~�Te*�E��Y��q��*Q�<7��^h�&@
D��S�+
s��S��w�O��%0�dM	o' �`�/\�^�$\�-O��=���$]\l��䃣]�5딊у��OD��d�.U���ݬ3#�`9¢
=D�!�d��\\b��U� t���!�$̻y�Q�/���F��Dn��B�!�$�5'Î�2�'
�0�r�p�F^<�!�ȹ4����N�"D�\\�gR�	��y��?�l����Idræ4O�l�O����'J�5·��puXY3f w�!�� �����0��̨!��1�=�1"Ot�*5/Նo��H��[�10\ps�"O��b�9Ldd�;GdӧL�p��"O�9(�']5qH��項��6���"OE�v�	�p��dJWET1"��eac�ퟘD���K�8��I�$�������'6azB)s�PC1�;5�Yi�)�$�y��ƺ"��a02�N�A�Ơ2����y�3e��ʂ*�`��w/U��yR"N�"�D�Agҵ'���#K��y�
KT��<*�̉!�|dx�&�3�y��9	T@�@p)�>ER�%ѵ�䓊hO����PR�ǉ+>Bl��c2i���R�<���5^��[���Vi�XIg�i�<��$d5�R`a��XFdl�6��c�<9������$">Za�\q�'`�<�e�"��1QSF�=iz~��!-_G�<�"*��C|m��k��U�!��B_F�<a�(L8�tV(L��L�Z��C�	3zF�q�$�c9����,��C�I�W32a�Cn4 y�xӇ�ɯ5�C�	?)F���`R:p8�H�I�}ffB�	�K����ǀM���c�@>DڊC��0-O.h�5l��uTܵʢ�	"�dC��9�b�X�e�9��5�D�˒ApB�	kЂ�@��Rn��(�;M���=���?���� � �Q��+/�����L�N�!�dJ
t���g%�B�,�%�[[�!�_x
���A&�d����1P"�yR�	>g��E`�9jL��%��,\B�ɏ/\���ɑ�o%H���-�$<�<C�ɒz��
@Ŷ/����hE$c��B�I�O���7��j��	I���3otv�=	(On"|zS �+z(���б1OtxrI@�<Y2/\-z.tc��
2puT$+�e�T�<aU�'S�Ɲ*!o.nd��;�d�Tx�8��t�q������Hg�h
GN����a"O�%��]/N���)��,��,��"O�-
��5��QB�N�q�R��"Ob���'4W��a��+�8p�q��i�O+��{�&��uL4��gR׸غM>�I01�U-T�dđ��!#>�ņ�/�t�'cQ!>�[��˄�����b�.>Є f϶V��0 ,]�z�ń�[!Fq�V-�
q�X�`�@�;�Ąȓ>K�ݚ��O�hD�����l�ȓl�TIK��� ����1"
�@GTDB��*~S�ڳ�V1t�� ��Ol��D��|�X�#lԮ|�b a#���R�'�iѥ��$iKT��!k6[(Iр"O��JƅւQq�x�*��|Y8)i�"O�]k�&��t�25J��ٱ~]�r�"O�}��H�@�a	d��w�>�K�"O�����>O�9�pR���T�"Oڭ���HF���W�ZaB���'f"�'�&ܐgؽH�8 [7D�}|z��y���)��RF�=�-	���P�?��'��<c�b0w�m�f G�s?�E"�'�pcQ*w�.4�V�+ ��p{�'(mj�F ^@4xVV*��'L�ⱠL�Ltni"��4Y��'z:��ύ
y���i��{ v%��'��M�0����Q��� A�����?��M�/�&ċ��7O�x�A�mK8�?���� �`2����X�h�G�X�h�"O`���&M�����5-��"�r}�#"O� F�ZW&�Z�k�0b�<-��"O|9��B�7Ɗ���*��8�(H�""O���7�Ϯf���W�ј!���T"O�I�՟?��9�'ŽB��3a"O� ���GQR�W!E/m�v͚&"Ot1w���N�9�鞞P�q��"OH�@��[�T���SjT�~E�t��"O��[��ˇ4,��Ĉb;�=x"O\ r-پB���Q6�$2�t �`"Oΰ�/��	N����%\.?��1 "O-�����X�����w�~�"�"O�3�,�9Fr2�S�3I����3"O��X�ne_��,�%,R�E(b�,D�ȸ��ǨbL�u��N�6��T��.7D�@��ۊ/H���"Ϗ�`���3D������&�r�#�&��\:1q�`$D�`XE�K�yкI��	�3YA6� �>D���茝G��`��K`�4yc<D���j���\��q�F>jm��zr�:D�  �0�F�(�K��9*d$��%D�$�ƬG%�V�v�C<�PH�g7D��yS�=[P\\��˜>K����d�5D����� ��@C���I�:�b�1D�(����?��𒔫�*�����0D�T# !G�M��`u�҇:�d��2D���և1%_H �ۅ@�ٱ��/D�Dz�ˏYk��RuD��W}m��(D�4��	�?j\��W�a��J��%D���q�^�T�R}�㨑>Id�1d�%D���6MU�7��$���f��V+%D�E�֤[��c� ����t9c�=D�����m ���5AH<�#r;D��qD�+/���%�!�<�&��O��=E����UQЌ�R�J&P�$�J�Đ{�!��K45��aB[X��h�`���v�!��αe��8��B���<$��:V!��gt��Y�I�\t��wBٴHM!�&b��W&$VM����I!�$@ȀB^�h�*) �]#C#!��)%}��@�a�r����~!�D�x���DI'J��H�gm��A!�8'�0�!t�	�"��u@L�(�!���X��h�G���-�!K�<`�!򄌪Z���Ru��~͈�ϙ�!��=�2B���46޴%ASĊo�!�$�S���(2��r��@ꆬho!�d�y�j���"̯nNNx(���,�"�)�FƤ�L�u����@O��C>4�J�'Xzp���8�@p�P���9�J��'�� ؔ��n3��"��CF/�e�'P�DC2O�����>a�|��'�9c��-N!����#;T�8�'���ys���6}����+]���'%>\Q�f��e���s�B [q4��.O�=E�T�E�	�4Ux��;f�p�Sو�y��SofT�"�� fE�"���y�A3�T9��IZ�s�Vl3�MX8��?��'3�<��O[�o}h@X�I���l����?��1s�a[�������=<�X� 2D��Sv	�,{"y���C�TP�R$%D��X�(ԔPfd��F��DP�z��$D�lrvˑN�dx����.:Ir���"D�� ,���$c5� �F���~���V"O~]��i�#�$�Yׅ�M������'�2J\�FH U 5�
�i����!F�����'�a~r�X���őG�
�n�da���y�C�m*A#�N�Y�Լ���U��y�ӊ`��D���@�I�4�5A�y��O�3	5���UGl��ٱgB�y��E
s��C1��A�ȅ��Z�yr�O��(!Z���Na\x�Я����x2$�m	�S�- w�B��`�I&���d��T�t��X���;�S�:�E�0D��p��K8
x�(3+�$����.D�tI�J u��%a����,U��y�C(D��*��˅i�T�e�
�e���R�'D�`Ua
�x:��"<E�p[�A D����E��j|���;Y�䑰.=�O\牐��e��X.ax�u�w`ʐ52�C䉺g�ų�N�e��1�b��;��C�	N�`���f�[PR�!�#�@��C�-[ D�w�ןs:Q
Ӫ�;���-�4�BeW=)4��b��"���c$�7D�؈&a0-��0�7�A�|��AQ�d3D�X���P� !���l]�s@�.D�ěc,^���]5���3`..<Ol#<������e g�2z�����T�<�8��t#&�߬uu�<�i�zh<��ҾgN`���
V3V�6%���S��?��0?)�lW/�bXh��)��$��IJq�<q�K�-5���3 ,W$���v�<yJ�� �V�i�C�fބ���y�<)��4(H�36�H�AB�(;�fv�'IB��G��L��@��|�04˶@�	^��B�	 X?@rc�H.6O�-ӧ�� c�B�[��Sԫ�9t����!�B�ɔN�P�r��Դ"�љ6�� �~B�	#<�f��F
�r�B�iv ;�C�ɜ=H��*^u��}9d#�>�rC�I�}�����d�/%��Re��Z$�?Q����P�`�n٘0�P���������"OXlPp�P!����g��w��c"O�قU��$�=sw���[\:8��"OBA����@��x�3ȗt�����"O�@ْ+!6�,�A�,@-���5"O|P����X���p�-��w(�
�"O40��+{�=�˃�j9���"Oθ@��b�cB��$
~��f"O6����R�J́�EQS/"|#W"O�-��ܹ�
+7���*����"O(xr`��%�#R%ϥo��f"Op-i��	��H��6�¸f�����"O�R6�ʕp}���/ݤb�4���"O��ԡ���| GI�:�@"O�xR�&�6|�jD���Ń{B����"LO��k��Q�O�0�:҆�	]�hq�T"OXy�ǣG �t� ��|?�L��"ON�"�b�)�f��T��Ihh+p"O�����~��uӂ�ڴ0�C"O��{'G%uה8:U�K�>����"O�"�E�:���0,N�;~U8�"ON�k�C�T��q��@����.�yb,��F�y�d��"���y",+<dD�)�#@�p/R��g Ӿ�y2��&�����@�g�x��R�yBU+O�K�D�'�`!�@��y
� ����/b�}�"́u�f!˅"O��1mO2Po�����D�Mڸ=��"O�m�Rn�<�p����B�t�s�"O�����[N�hP��iB�5���p�"O���Ő�ok�`!�HB,]��'"O�E�w�Q(���፠I
��"OVYC *L��9��V�V���U"Ox����?+�6�(�۬v����$"O4���ge�<�p�e^%.�8�3"Oe)�,B���'�߹#kv�!�"O�XRG+��p�d)R1-��@$"O��	��yh�`g��7~@T"O�ⷩY4M�`A�7i,��k@"OD�r�0�^RVH���Ыp"O�lڒ�Y�������E�[��y��"O�E�pƷCh4Q	���R�>|��"O��2�&M>�
�x�O��.nZ��f�|��)�ӳ{�$m��䙫B���y, 	C�C䉻G�@����
@i�q���MxZB�1��v���� '�"46B�� M�^�QmT�je��р� ��C�I�>�U3��^��C0	�=ʄC�S�:�Bg��Yw��8�~�����	�.!,a�I]玔 �@�YzB��.¬�摖/o\��f�X�B�ɋr�|`��N�	jKJ�b�<9�BC�	� ��h��"�@�9sF&a�2C䉝KWn\a�)�m5�$*��:�6C�I�b�0$ir�-�X4f���i��C䉐I12�Qb�]�# H�z�c���`�?�����n�&ۤb���!�+�6[0!�$U ���RA28�x emΞM�!�ыdx��# �[�ٛ��D9;�!��7X�&u���J��`z����i�!��
> �2ɖ�}�-".��w�!���JغDE�
hn@sg�\�!�D
�iF�̓�N ��aK�>F���q�k��~rcٕVd��M9o��r
0�y2mU�W��0t���V�L3᫆�yB��*?�z��r#II#J�0o�>�y��C��j�:P)̞=ĐP����y"$�1A[,���5��%�' 8�yүK�� B¢>!�99�Hڨ�y�,�.��SGiX�*�𔱦�����$8�S�Oޑ���։lp`W�]��	"O*}٠ 	S".m�a���)p�Z�"Op8���8b/F��t-I�AP"O�P�v+�0C�­����X��M�"O�	����)���RD�`�����"O��q�A1R����gL"��:"O�)pd�W�I�N��� %�D���|rY���S�JJn��c�7R hy�@N��H{�B�(t���d��M6M2���k�B��0��H��Y�X�A��NPu|B�,>^q�D^d9p��7y&C�ɦ�誴��x"=�� I4(_C�	b�"ac���b2}5-߸C䉣H�t(���V�,@���CP
7K�B�/���!lS9'r�Չ%:��B�	�]�y��-�	*@� ���t��B�	�L��p���"^�^�
C#Е[��C�	�6��%Id���-]Lh�2
�tB䉽2��	����:.z: 0�����4V���É�V�FH�#�]!|!�� dŉ�iݜ>�dd��mU�y���r$"OrH ��Ԍ9Uꐉ�E����
�'�'�B��~F	�y�ie���_T8�����V�<ѵ%�)�\��NL�ʕp���y�<����nd�<j��� �|(�)Iw�<�cD��,�����ps�л��[~�<!��:dc8��揁!��4��eS�<I�R$�C��6����MLh<�*��X^�I�Ce�(ۂ���?������hO�I��-��a��s��� CB�V�!��*��Ò��j�|"�"Be�!�D������훴4|�h����*�!�Ьв���'8~\�����_�!�d��z1T@�gK�|P~܋���[�!��&/����Jް~4�z�ᝒ�!�$n��d�� Y'���Sㅽ��Ih��T !m��Q�h�@��A�o�L	g<Orq�Bቨb�&��!�[T���m��uY�C�ɉM��u �E��e>E��S�@W�B�ɠ 7i�2�)g<&Q�u���*C䉈eF�B0Ot3��r�N�*KC剮,3�*`��%p�L���w!�dд'@!�>X����ć�x�!�d�V�VEB"�L��X�R��t��y"�	�vvJ��%@]�ڹ)BIePC�I e}��z���Ⱥ���ާGt�B�ɮ^�6d�.�v���)S偁j)�B�	<�*-���l(��j�ˋi\FC�.y�t��@�v"�H���ThC�	�{ަѱ%�)'�,�I�FU�_3<C��Uo2L�T��8Xj,񓢑�!�&���W k/B�!3O֡�-�+�HЩ�Ҡ�X�"O�9#)��s����eDs&�R�"OD)����r.�#Zn��"OlUy�CZ�� � M]�*�x g"O��	���1C����l2,Ѣ�"O��ٴ%�Bv�K�
.D�}�4"O��S5���d$Bh���5�;���$�����x+�j��z�'Y��xCUhH'6\sw���~�1��J�[���
9#y0�PÑ8;��P�ȓ9��4�.o*�K4��1s%�����D�O�Y�r�{D�^	d����e��p�(
�|� ك ֆ1�I�ȓiL< �!G�3�UZ H�X2�9�ȓZ�|%�@�S��z�p������ȓмM��ܴ&���W@ƶ<�݆ȓG98X�E-�y��K�2�NɆ�X�R]<	��h�$�Ŷ+@0�ȓ4�ν�/�o�Z�"s�=G�F��ȓB
z���N�1�׀P#Q��	�ȓ.7^�&�Ѧa-���4���Y����ȓL`:!õ'o`1KtCҀf�T��'��{���8\8�]{�@D�I��q�ȓ`���#̆#ɪaad�T�T��ȓ=0��j���m�e��K)�r���5�i���1uj!��8u8�����z����c��MhCe�cLrA�� ���*����T{2ȸ��wh
e��9���3�c�������@�0�T���	(�IS��P)������+� ��pQH����+"����B�|�@��m� ��Xt HQ�Iڅt����ȓeBX0�S��Huc�R�2F̆��X���˕-7`�cVE�Rl1��S�? �����*]^�᷌�OL�M2F"OR�9�D@�m���y�,J@���5"O\��^�q��Ԓr˚	$�
\"O�}����&-kѠ�+�b����"O�	pC^��)�RjA�l��"O*9ڐ�C))>PQ+cH7ZEi�1"O�M�$�9/�%CwENg����"OR�PT�ǓN��\�G���[�Dؑ�"O����ԧv�R�;b�X�H��"O@��¯3Z|f���Br���"O�p���
@��k���a"O�����:%� 0vM��f�@Y�E"OtKQ
hpjW�Ը2-lDc"Ov)�%+�pj���T�����1"OJ�k1&Ċ:�!�d ״B�R�c"O��` ��>9��H��@�.�|��"O����s�~�jsb�&	��t"Op-qe�Ϣm'lqZ����=��""O�y���m��)�O<�,��e"OD`��&R�1L	�k	�{�T��"O�Ūd�̷+ulM�
f�~�0$"O�)�'F[�[m��1���"�&|��"O�Dl�?3�i�&FץM�� �e"O���Q��%�T�AЦ<�>-s�"O���F[C�`����(	~T�W"O<e���M�F���C[�#��(�"O�H;�OI*)�[�B�0��"O�dh5 �?T���eU�p����"O:})AG'�R0FAqP�C"O5:H�4c�P�&#K�*���;�"O�5��aۊN��@��b�@�M3�"O	త�[g�d��@��r�KQ"Oh��v���*Ap�/����e"O���l�<]-HhZen�#Z�R�"O��q��U/��1N1zL@P�"Op�r�����)��ɥ8��s"O8A�^�;m��ȱ���F�2�`0"O6P.[�v A��*\���]*�"Ov�◎�8t!uP7d\Id�q4"O��Ԯ��* ���Q	��\I�iy�"O�� r��:���;2/�+ :�-�!"O҅�sBM�cHd� �N+���"OH�	f��n�,	'��x�NlB�"O����=<4���$��D�"O4x���-$�Q�D턨+��58�"O�m`0d��?2�Ő�k[	̸�yS"Oܕ�HZ�Q،h;'�ޛ2��r�"O|���DҘ �y��A�)���ru"O�!�Lƌz�`MPݥ0�d"O�	����U��8P�� xi&aJ�"O4hp�)T+\���0嗩BE��11"O��ӧ�VS�8 5$��=L��P"Oܨ!LL�#y<��W���^���"O&5��ăYGi"uGU�9
J�U"O���G�24��Y�v�0�`48�"O�����,Ip�*4�Y�z����"O��4
Z�7���4��
aTh3"OF q�K�v͌�z�o�L��0p�"O��GA�0��,z�ml��aJ"OHY��&<[p!R�M��z��i�"O�M�S
�!wL� �ҥ D^�bW"O��W�@*��P�E:��ّ"OJY %�ʎGw�����{92���"O���̽S�z�[s.�*sU��ۡ"O� �؃�ژ�Ny��.:���"O>�����8`�-J/�(�(�"O.��b��(h�A���0a�|R�"O00 �M�(!�����?$XN*�"Oz�qCZ�Z����u(	 .�@�*v"Ov9��G�&�2h�B�0`}��"OX�C3��7$mہ�]�6�=D�1ǴC:�5��N�{���*7D��9����k:6}
��5�\<K��5D��a&�6�Rp�0H�:�btA2D�P�P◷�x�1�ڱ2�L�b#o/D� !��D0��<�rT#O$� ���-D���҂�$=��;�/�?���Q�i'D����I���`�.\��d�A�%D��
N0��aCK�&Wʴɖ�)D��J�����B��ψ�,N�p:D�d�
H�Z7H,Sa*�B��5aG9D�P�փC�zu>e���Ç�%��G)D���-g�& �Aa�6	xA2D���� �M��̚J�P��q�=D��q'S����ˤF��l:D�8��̀\��}2�ɉH��H7,9D��ٷ�0��X����g�����j#D�@�"�̗p�;�hL�X:mQ��#D� "��� 4Z�H��Vvg&͘V�?D�h�O�v�B��S�X,Ш��K8D�P�P�C�[�>�;���	��M�55D�а�
�X���͎>����a�3D�,�D8X�Y�������;U�%D�X"U��&�"�餭T�Z	�9�#D���E�0�t�bS���PC�g"D���`�_>Pi����Gp�4腋?D�(��$H3�X�ϐ�c j�5*O0����ԢV���P��"z�$Xِ"O�ݚ�`ݼu�m�p�*
�� ��"Od-��唬��񹕡��}I𔘑"O�y#���"�B��A 6
�3"O����_����HEn�!�����"O���6+�0L��1��-{��a"OT �df�!.�M����?f�"O~��F]v�R=ڰL؛"�r�y�"O���m��T<�N��e�f��t"O�5B�L����F�#\�.�!"O�	�'mE" �|��F@նG�0u"O")��e``�$�U�c�n���"O^��� ��+�
%����-���a"O��qsM��%:�-`�KQ�0	�3F"Odh�.&�3�H��4e�T"O�k�00;rQ�eIJi�"Oɐ,�b��Y�ܢ3+�X��"O  U)҆"T��y��_^h�a"O�yv)ܔ��(�����!v�C"O���&�G�օ��i�hY8��"O��bP��$rDi�HCLJ4��"OD(1�me�J4�&z����L�<����Ho� +@���p%5�Aq�<����V�X�&�Q�,�04`KB�<)B�0fO���n���T�@Μz�<��C����;�M�5�0!�U�s�<��J�(Ť墱�C�6��\�%$ x�<��%�	ZĲ��5,�$|����#�Z�<y�(p�jt�E#[���Yԣ�y�<������H'���.����o�<!��+�@T+�+�$Y$-:���S�<� $t[���H|`C@ƿw�
���"OT�SI�
xQ�M��؞8ث�"Om�BLI).���:D/э]�:B*O�Lx5G�Q�TT����t�#�'��`�pB2#܀��" ��	�'� @E�N�|C��
'M�]�R�'0��`� �N�3���< �����'�@�au���땏��n�ȑ	�''���p�E�ƈie���X�:�S�'��uK"��{�	ٰlS�_�T��ȓDt"DcVŬC4P-u�!JG������ha���9�*�i�m������syJ��$Ɗ)*��1�nS���ȓB��r��ݰUQΐ�T��}&��ȓ@��,㊊Q��D�C�P#�͇�t|�]�f�մZ`A�v�YZ܁h�'�H���#~:�i5o��h(�P�'��Tx�Q�R �&T羱� ��e�<yCa��d�B3b��"`o5âmH�<��J��=s�%��OK�dKj���J�\�<AG�I<r~N!���R�b��e9`Z�<r��*c�ڜ�T�I"-nd�Op�<A���75��9W�N�(pm T�L��헒,�$��cJK2�.؁��>D��QF�RhvI���)L���1j=D�H���HU^ �����? l½�a�?D��K#��.Z�<�;֠��k��q�w�?D�PـFȺ| \���Ec��K�n9D����''��x ��*�$D��)''J�(þ�ɟ[U�|�h.D��F�Ҝ6�D��e�'o����4L0D�䡆 ܵ#��UA�Bx�����!D��B�3@�M��K�=Va�Ԛ0�>D�|��I��?P(%��J	9���c`�6D�� �"'*�9íŎ!�
�_B�	�$�ܬ����)Z���o#JC�	�/�攒Ӏ�x��h�L�af6C��
U���Vh\4g�z��P���+D���1˂��U@��ж=���)ӎ"D�t�PϠל�`B[�2��)yB�-D����g�~d&�*������u�,D�T���$G�Y�r��^�����J,D���TJ�#7PB�4!���")D��G�=� ��	`t���`#D�<rr�C�`�fš�#�2¾���"D���� �kvEJ��2s(�)#`g?D�D����C�|TA��U�	' �ڳE D�`�$(Ѯn��� u��b��{��>D��_WӀ('�o�z}�E8D�hY��CP �$��N�Z�B M6D�`�O�J�� y��<o�HQQD�5D�,���ӂ|�@��۞R_��pe/D��9��'j�5"���ӗ�9D�� TT�w��y)��3�h�@!7D������9��;�l�#(���5D��A��-��a�e��+[hJ�(2D�\����x�u�tƊ�ls��jl0D�*���#A*��{����G/D��#��d?��7Y*3���s��0D��@�e�&&��Ri�>RI�E�n4D��2vI��p�2�����M�>D���B$�:i�
��ՊO�BU��ti?D����Z8SxR-�p���i��H�>D�(��)��9��Q�`@Ɨl��0N;D�� |`bLw9�U���4 
>R"OPD���)�<��@���?��Ij�"Op�P�b��eW�tq$I���9��"Oj0gk\)� Pks��7��Y� "O�i$N�8�i&�Ƞ��c�"O�[��*˪L��/$
¬Ī�"O
��RÑQ�TYp��ܫ`�"M�t"O�|{�N�q�p����j�l�p�"O�(��wLHؐ`�("�Rm�$"OD�Y��7�pr��R�Nx���U"Of(J�-E�ZMA'�H�^^�m�"O�5��G�M��&����  �"O��c����p�pEΦs����"O.M�!��;3���q�۞:��� �"O\�{WD�B9�%Dy�Q"O�U;�n����@$�?UkȈ0e"OX �*����ˁNL�A#V"O�M��ҐE�\��@�I ZK�:�"O�Zq%I�{�и����\�(���"O.�I�GF!B��4��ȉ R"OڠX��QQPD0��%V�R��U"OL�	��K�Ƞ��LR.�豠"OF�ru�0jX��ZDf� �֨�"O|�3���)r,e9&+˳�\�ȇ"O���'@��L�Y�u��(�>�A�"O�5�`/J�-�Xī� �Yf{�"O�mZ��'Z��^$���"Ox q���658��A�;)�Lu8�"O4��SX�bR-�Ɓ7SB��!b"O$� Q��{Z�1FI�V7�q26"O�����z�R� 6Q�9��u"O�����[̒8�����Tِ�"OJ)	��7IE�!��c	Y^mz�"O& �@nן.���B���Z�"O��0�H�8"��fX�>��m0�'�ў"~jt��5c�BdA��1��R�GB�yr@�k�
A�\*.���X��ԭ��?��'��xa׫D�mL�l�r�G���'-$����	.�V��p��:<}��'~�X��i#	Q�}[���@ʹf�!D�<U�߶uz4���k����g?,O��<i�ԩi��L
���	 �9���}�<q�>L�8LDy!����iE|��hO�O���'�e=Ja22�&k�\�N>I�Q
�,�/R�M
�X��X�X�R���Bx�۠o�-+�4H{$Ɖ�l���ݶ�B%��*Xu�	׳<�8���ɳ��'���)��@6�����M�b�zy��'i̬�i���9��@]=`�.��O��ɚژ�H��-�&R7A��X
��Ţ!���j�"O4�IƮ��z�����>0��hr�>i��O(���
4S���.7T;��T�Q��E|��O8��WG�N�"��wN9F�b���O|��]9F�:��� 8y�r邇J'��x��J;Zġ0�Mp��������yb"͠[�%Ӆ旛w��QQ���9�S�Omm�ʏ+�$�7��b����'/L��M >s'�v�� �7�y�A?Uޚ�ٴ��c����֯Y��y"��
Nw\�Q�dΐT� �0�@'�x��N�d��.�Jr&�`�b\�=l�
�'����	۩?_��0��0Z"�5�
���'�z9ɔ�L7zV��F�ڏ\�x$(?�����>V���b�^.OP�)p����(A�A��⟄D�� ج�G��8�V��bǐS̱�"O�yTd�(Q�a�,�.��yC�It��{��۝*ݼC�cͽ?�ɂu��[iab�O �JehO�>�(*7�F>$�D��'����ڲ)]�5,NL�E�֚X=�m�(D�� ӈ�R�
���$���kF�0D�;�B\�h�p��/Ô2��i
��!D���'FT�5���ɰ�$�A2�b=D�D��$Ė�B�%��SB*���<��B���t�'~�n�)O�������cbҠh���d�a+ܭ(%'A�|��J����X���hO>%�����+HD2����9?��2tO����2"r(�Q`\.�*dc !/��u�����F��Nghg�ZJ$x�5�,<O���dy2�i�4Xawj�2WWN0��Y]�;
�'E��+a��xC�̒���!L�N�*Oj�'[ў�'h��a�%_�j�����D�[����G���Aa�ϛP��a+.j�t�O��=��r\B���` �G�hx�e!�y�<����?k�xCƊ���d̗��'�azҍ�]=�c�	
�j�3uEʘ�y��#��Ao ����T��y��A#F��%�p.��ژ�HOң=�Oqf,sDb_
C��I��/�⭊	�'2�B2G�G^ɱ� !s� [�4�hO?7-D#~~b�{���5�xmRAn#�ab�O.1�"���S�f���>E	E"O�X+E*>:h�)ae��ZӮ���"O�,yUfJte"`:�Æ)'�isüi¡��E�`��Z5��H001K!L�%V�6�)���{0Ğ�2�N�yt�8�b)(D������/9t`sg$�7���֭'D�Xy!bT�B�,��Lٝ�����'D��[����$?�YA�(L*J���k&D�SL�.P��	��9�E�1D�Xj���>�(�4A�-�j�*/D�P��
�,�T����&WCF�+��hO���}�����5LtD⣈�
(�B���|�����0�6��$$D���6�g?N��	�˖�P쉻� Tl�<����N]���t!��<�K׎��-�d�'F��6֙bxD��/�9�I��}�A�_x�����J3o�l��	��Vj�ڢ!D��
���	*n�I�P�W��sqh$D����B"f4��P	/T�x	e!D����� �W��s�o�'RJL	���$D�,�dHV@�8ɶ���$p)a`#?D��&�ϪcV 	i$�l?�4G�1D��Ȇ�M(Is�a[� Q��Ȁ�D1D��Sge�0��-: M�ƴy�/.D��9��_�K��I��1���G$'D��ہf@�}J|� ��w���&D�`�� *\�U�Ba��8w�`��%�IC��tqmяb"xU �.ZBZT�/D�����p��[C�&t+&@sՠ-D�Ԫ�!�]�$Y���S�@��yA��-D��B�IZ�H) ��d��0�[�&7D�|JF�W�O�(8a��4H;��طȴ>	GA�KX��Z�dp��*�hثh�f� 1�2�OnͣRT����)��>�U�7�/ϔ)�ǰ������o�
ȊQm��|��	iSC�9����d'�->7 Mr��I�WS�}��[�IU�B�I��촓2n0[ �8i�	�+D�p"=	:�I{��paq.J w�
}xf�M3,i�0���� ذ�:17����Qh����x��)��$0�x7�L�6�<qR�AU�	>FC�	�P�:��",l�"d,�Z��7M(�ķ<�|&�d�3�ݦShՊ�Z27��a�<D����͖�	�	Hpʗ�w�>tZ��>���8�2�kC	�E;�i��y� t�ȓpG8���N@:��Qe�i�ȓE@:��s�E	-Q��v��.���hO�>ţU�M�@��arQ.�|Jf����?D�0�&LHM7zܺ��7J��	)��>}��'5�����;Ƅ}ː A�{>$���'vU!My����H�w�T(��'�$��d�$>q�P��?DH��B����zӞ�/�p JEʀ�v���#��P Ԣ����nT��K�>[ �T�1����Dxr�)
�� �&lX���a],���+�C�<a�O�rh�jDkԊ'X6���Ju�<��ȕ3J�"�J��V�J"J(����w�<0DW�vPڕKu�ozZ qu!�p�<Q��=<!��⮗ �>XB#�G�'�Q?-�1�c���q��?p���#D��*rGX.6�\}Ǆ��:�au�>���铫_1��9� W:j,؄m�$'"C䉮+���aO��Db�G�#o��C�ɓ�`\KV�* ��4���M��C�Ɉr��A���S���z���(mb*C䉟_~޵��X9}Gh�Ȥ&�4N����d�<4���v�p��� q�"0�B��_�<�G��6�
��S+�W��8�FLI]~|��8s��᱑�O$SO��@Ƶ	Y�C�I7��� �IƇ[�`�KE�U��C�ɐg���A�L�bh���AjL�C�	1*A�x��)�,ǈ��c�$�8B�I+6��	Ce��rl���<q�DC�I�+��l�b�!�L���g;pC�I=ldnd��Eʅ	$X��o�K�B�I�I�;6�d
�Ȕ͌0n˦B�h�N% ��h�������"�B�ɎMR�����ih�@[�HB�	
M=xTE%ԝf@ ��@"F�4B���Q7iը�,�0T� }rB�	;����`�VN����k��5��B�	�J����j�H���>\��B䉵L.�����7Zr�,9�L �Kv�B��7v"qH0��*<��%r�+ =-�<B�	`�
�HP�]#R���
@AR**B�I�IHa��'@b|9�gB�+�B�I�g;������-��H�RB�	�1�4��CT�.�,���.���fB��,��}CW� 3Kĭ{7n�9_R�C�	/_\@4���X�_=ĭ�J��D��B�	�KGʽQP�Ą}� ���_K�rB�=���%j07�}Z�e�bg:B�Ɏ3�xAB��_ J�0ms#�B#yB��%T���h��*qv	�D�ޡ�B�IO�z�q�K�2r.�;�^�K��C�`�� Kš�/H���ɰ[!>G�C�-18 85	<D ��������zC�	9��J��΃x�PXk���=i1lC�	 t�%���$R��֧�5�XC�	s֑�0J�0#���b�Р?�B�I#K��`�o�*2��Kίt�C�	�P2
x
wA'M�.)g��&��#>9㪇�H�0T�Ti�"��ii3��<�5�G�*s�
�-�'t\h����t�<� �����V�%R���2�|t("O�e��ͳK���Tn�*@Ґig"OȈ( �,%&1:��?�xjU"O�J۵w�(�m8�Z���"OF<@"ʄ>R2b�q��V09�40 �"O�$�@�\�F �IF!�c�ěv"O�|Р�^�m���Dc�84� R$"O�͠'D�(�d1��߷g�L)�"Op���&��Sϒ��g�Υ>�4,@Q"O�	�a �l0��C�9~�%[0"O,T����L9]��(��`D��e"O"к5��9r>={1�O�u!εв"O��J�L��xm��ٲ��Qp"O�Hq��HN���\wlxb�"O�i�T�d5�U"C�t�.���"OH�+�����	aBC��6�*�"O��+�D`;�CW�� �z�)"O�!`0��[�����Y)�b��"O�-�A�#+�>���_��&`��"OD�:b�@�fp��aE�ּ��9C!"OF��d@C�*�(�ǋM�b=n\�"O�̑�h\t6���hX(�t��"O�I�� ӂ�^�h����_�ı�"O���^�; �$"C�H*.7NR*Oڭ�������uc�7�
�'�Y�b
�o7h8J%�^�o����'ǂ���O�5p���re�޳o(�<��'n�Qz��Q�NP�4�F+���
�'>��į�$I�9�'��[22�	�'*��xca���:�p���68�
�'D2�J��S��i�L�Sj��S	�'�r-!�E�ZVN��$�GLa���'�ѫ�,\�+��Ui�I�x�
�'��z6��@Z4����W��'alH�i�=��j��TR�'䦭X J՝B�ZT�7)��
T��'� m��/C:F�;&JRh���'�R�p���<;8	�EnT�z�
`�'��}��,\�J,+e*W�J�bъ�'�6��7�D��'r��k�S��!�߆'�\Q
�6;��󥃟;s!���ay��K��B�ij@�C�9S!�ǽ$YR��ڢ^���o٠:<!򄀪+Ђ3�Ƈ_�~e��/�r!�#!��(Q��'��ڑ�:u!�DZPH0��(Q�`�P�+�*t�!�U�Zd����b����Wg�!��4�
0��߅R���I���!�䀐@��mjF�Mt�����I�'u���Ν�H�xҧR��>�1�mV�UJ��	�~؟d�G$d��y�,]F����<\^�4+7m��6��b�L0z�F���.�4�J��^"G}bfX<b���@�Gl$�O���)v��7�B:�χZ����'�M� �6�ZRM^l ����'�� ��V�o�2x#�W��}��'����ƀɡH��}s"�a�<���PR<�=�K�1B��	X0H�剬K��
 �%e��g��W���b䏎s�f̒S��-?v�Ն��:�d��DH�Z��IEb�m��9��� �K�n��U�Οհ?��̇�`U� d�W����Dh�'�� ��C�>^Y*8I�du��#G�d�r�����55���`Ø2��tR�
O�Y%���G{�h��)^&yf�xC�'��8G�.��M���76�A�E|�t�ҙ�$��q]�b Ì�\�����t�!�*�z��l��$h�ڔ��$�ޭr�Mǽ,�h�C bV+H�Qp�Y>%�U�
\�.U�'�&�hwj�ƈ�D�gb�A��fg�i���S��� ����m�V���@ɘpSXg��0YH�Ɇ-D�\
��1���v�ax�E�+h�����8o��%�Z�hO�h)T�[�a�M q�{Ӛy9�MȚ-�Pi�D�],%�j�)�30/N���CM>�Ɇ�,�.�س�;W�*������ɍ?:��х�VP�l�>R�u��'�u7��!L~��K��!���a�	l>�)v$�~2��QHhS�Iq���)�� 	֔T'׈W���+ �y�x�:PA��r�����W�q �=�Oj��㫄*]\���l�R-��#�5"p
�14��:�
5�O�����=������ {f���*Kf5 ���y�ְ~H�$Q���ѥ� 9�G�p?�� ��%�D8��W((��6�	���AR
�A�|�,�"2�Y��%��e޼u�<}�˓-'����e
Z	]��Sߴ��'l,|%�|2,�+s�U�Gh43ց��
-�O��b�i�6]���C[4��p�e�br����P;y<:�Ѕ#[!T^x�a',O�l0#����
��PA#��O�d,	�ap�� 8$�O��8r�M�,�]ro��S����5�̇"!l�O����j �\!�����U!���<O���� 
N�|A5�y����A��Y&��~����}iZUz�l�63�eP$A�<9f�ĦRu(Q�s��>9�eQ�a\Dz���7=XА��ac]=�Op��q�#�$u}�ո�j�|���@�$C�a~B�R }M昻_Y�����$��K�.mK'd\�v7�͘���.XI<��R7v@���ơur��vn ���ό������\�ڱ+$cշc������A��4H�,�dN���F�UآGCh<��  L:�t�3�ռ�T����F�<��M�=J�Kae���,
�	Є�g�OV}�%\"Ti���d�"�'�]"Gn��K�8Җ�g��0�O($Y��A�Ȭ)�	ǓFv�=���O	;Ed<�0AG-/{Ƞ�?��%�u���?�1�ќp��h�A��m`�u�3K�-GI*Tk�G�VH<��T,(�8A�_.ҵ)'&;�JA�B.��ںuA��8$L��X�o�vi�S#��sw�M�-�B䉣j1����+V��.$��r�#j3�����T����D =NY���s.T�c����B�'z��z2m'�<�P�	��<�U��j�R ��Էsu��{�jRq�<��E�If�PSΆ/4�R���rܓ�f���X�������Hx�\�E!��m."Y!�Ζ�̐J@n�?SgQ�P�SX�\����(��-��|�'}:���1�ŉR�ֻ+TT��'f��S�.r_<8��Ђ4�r �89op�BW%S��?�!m�#+b#?	W��M#R����Ж�H���Q��pԥD�"v\PF�iv�DA�H�$�u�lǞT:�c�M�&��yaQ�'��0����s^^��E�}�&=!�{����X����7ǉ�0��Â��.o
��O�d�6�	�8�Z%B�G�q���P�'?����d��kVR���z�LQ���(/I��nڊ?�.�(���!ʑ>A�'������|CW�#C~R�i�'t��Z�fG�ڡI�,<����G�n�xVd�O@����P�����d_�qr醫1�2��v��>��DĮ{N�i6��.N��I�+�&E��Gdߛ`�����@� �p�ʳv��X�eO2Giz���I)������V�o���!X�%�s��0� �Z��ػI-�C�	�Q��ѰU/\W�Aîُ0���'��0b#�ܱg����S#X��:��� {��|t�O�dB䉡Y]:h�	���҂T`d� ���#}�EW�����}&��A�/Z4��@J#��(P@d�릭/$����D�� <9P�=�A��i�yN���O��<�� Z�����D۬B�1q'�G�WaXh��D ��y2�ǺVc\l�	!����d��H��0mӫgH��_�4�`AQ�O��3�
�.q�d�3��
>�Z`���2c�ʵ"��%[�Ju�җ�T�O R���!�}+�U1�J��y��Y_��(�Cģht�T�"e�8�M��KP#`r�PD-N�IZ�� ���ͥ,Pr���6^��h�C�Z��y�O�D��6\��ȥ�@���-c$HQ/j��Up�U?\\<SЯ2D��F�T�V���e �t�^%���:!4�JC҆hz�G�Dηh)��kM-I��9�SA,tK�-8R��rĉĕr#,D�˃�'�ڍ1�'L%!� ��I�d}*��?���y,O"!�u��*G� ��g�PN�C&S!]��ď"B��+o�,�C�ꍘ.o�d���Y^�<y�e�*!(B��A�H���8�"E[ �"�"�#�����F�4rL|�A	���	x��� ��ɧB�UY�$�w[4y?��q��'{���gBJ��F�*r�#Z X�PE� �@b�0�@딪 ����
S8XB��K�
�L�Fz%�����fO��!J���On��ƣљ;WNl��&�)5@�t!��d�*Qh�$#Ϧ���6M�@a1 G��|\*�L:�OBd �i��@��c�7� IC�Q��#��=�����T�a��9V��x�3A�H�R��1�Z��ᚑm����R��DB�	<Q���5˫O�p�%	� <v�����\I���D��]����W�Q��ʧ'�`Q�C(��y7H�)gy�H{wē&6��9� �x"��e���ߪ8�x�:Qj��.���c�ibz�{U�T-\�q�Dy 4��Wt�l�I *)Y*��Q�(M�����8O�l�Pƽ�0m:kK�f�RTJ J��5r������9��[���a��ǚ+ћ��'�����I�#��
�@_g,ѹ�{��'��L��ͶIH,P�eԁ~f����|��ǅ!4��d�w��T12��k^m�<�� מY*-��*6�˕�	�/	v��`�z�`�����^ʚ���^�i�|�]�|jV]A��Ƹh@�F�G��C�	��)x��+Z�
�QA �* ����b��F)ʀ�: ȝ�/��g�'�����?cR���K 2@H*Ǔ��$�#,�����7���a� �*6��{!�Ws.S+��'
����Ϫ]A��	%�:���ǭ�ў$+d� �h�L KA"I1NA�O�Ptz��ߪ`Ѱ��u��8riJ�
�'W�Iv#K�I�h���,��\��x��'X�D"w#��g�h�O�>q!�FW)#��ͱ��H1a�n̡Ɓ:D����f"qI���jӱS�^�q��.�D�1S�\�y˓[N�<8⎨VA��y�W8I2�`��]�A*e�]�_��)��5%E����3�����mF�A�y��W�	�(}��I�n2Q����iB$=YPL� ��=�x	�"n'D��X"�U�R�	��e�p�t9}��SR���OB.��ԂN�]~�+1Ú+}/��'�%�r�4A�1�U�+C0)zѩ�h�<���)Py2��ƃE(�l�g�i�����(�)+|0�2�3'	a%+یP��'� Z����I����I72Q*E*u�$���4p7F2ҧ�3���ud� �#[(P��H�ȓS�r�Y'���>�����'@/W��	u3�l�#��S7"��fL�;G
�a�Z<�Z�ȓ	�Ё��V�6�@�	U��BE�<)ČE�l���W!�X�3[M�<���ՁQ��ѣ�Z�2�i��@�<��j=|ɬ��ɓ%~ڍ Q�YA�<A��ԑ#� Y�g�'�`�r�Y�<d�� ^ܪb��9�ApW-h�<A&Í:�I���=:@n4��K�c�<qA��>���*��G5^�@Dz�,�^�<y�CW	
vּz3ҷ(�~���C�Z�<�0jر$N>m*&LL1�~4��A�W�<�$dY.S�jٙԡG�yn�y⤘N�<qQ�N��d E���$p�!��D�<��gӉX�h!�RD�]�`9FC�d�<i#(
+o���3ւVr�"9�'cz�<	��D�I�0�ئn��%��şt�<A`��C����+H �R��r�<�o��yR��(\��x���Ao�<��#"������w�l�" Ag�<1�b̋/���*ƪa��0��g�<���n��@�3ǅ�-�z��C�U�<�u#�(��͸V�uB� �N�<��Iw��nV�0�YH�#��yb��	�n܊��(7$$tRjҤ�yRI�$ܔ|�f���G�h��Ȧ�y��̪=����g�9J��!�b���y"��w���[5���,̅qC�D%�y2ȗT�Vl�S# �Z���E��y��"Z�2�H�\�k�4co��y
� )���"-8 +C��x[���c"O��t��p�pJ$ �8V�� t"O�Hs�/	3�$����@�%�T"O��ZD��_���F�*F��CB"Ol���K�P���@�=��"O�� �
H�X������'�>�9�"O:��Q�O�l��"�~HX6@�.�y��֓�	s�C���-�5,W%�yr+ٞ(V��&��.�=:U����yB��-J,�i'K+2�ŹD��y�L�	l����R�d�^�@�J��y��Jv�Ж����D�	�'�y�	�J��e���ϖ2�<d��	�y�e��D�$��T�9P KЉV��y�&�/DEt�"�.�H��`s����y��%����b��G�訒l���yB�^�-�`I�%�)`�Ȳ�S��y��U�#Q��j�k�����@C� �y2$[�CN��-�?�$0qw���yB�HxU:''��e��m`�g��y"H]0E��1�N�P��P�B���y�悹SҸ��E�N�$]	�J���yB@K쬘����A��!傯�y���j�"h��<=��p���yRdE���< ��1��P��4�y�� V�<Iǂ�6�� i%�M��yr��j�ⷣ
�"���c�)��y2Ϙ�}�������%"��V ߖ�y"��9d:����C$����J���y�ߢe�.�BH_�#��E���ё�y�@�&F�v�Ȇ��6/�i����y�H�
;���x��H
.��<��'D�y򍅮y���c���$�5�	�y��J0�H��2fU�S�����3�yBk�akF ˦�E��5*U'�yBA��9� ���Ȟ��P���P�y�`(Z�P�A@.T;:$�A)���y2�J%@�r+C�!�5�`��y��>�L��4�݉�R�c�ɞ
�y���2p�c�K!@�)���T��yr KncQ#C]��H)rc����y�n3� �v��b����e˙�yrgل;�N<d�.Hi�E�)�y��^�	k��B���l���Q&I8�y�`*:Mۀj]�0:ݲA���y��˩0w� �ͅZ��`��y2Œ�[s^�MLU-���A���y�	0"�x��ٸJ�0؄+���y"L�0R�P���� L:��cǨ�y�YiVT���W}��yq�1�yR��8\�Q'�ۅw�X3UnA��y��X;]������>|��̘Ԃ��y�NŔ��!��<j�.P����j�*X��G���0<ɂ+�/5<h�Q��>(�M1��}؟$�ץ=]���W@�(�൫�@�~E\HhGo��r�7 �b��5�HS����H>��Ojx�[�n��aT��ħT�>�zcBO�t� ���-ջ3�pi�ȓ%Ȧ(�n�7GN��¬��a����uW�"2�cM�+O�>!�Dחq���	�A_�y�v�K�h;D�C4�0b�6,h�h�_�N�)�!0����"r%d=Z�'���3��5Ƽh@��.�h�B5Q l�����6P�@��­j�&���E?��$��޸;�4��f̂|؟�1梌=>�<�����/&��"7�8�ba����8I"���� �)r&����+`i@f��+b�!�� 
l
�n\�ZA���'�H�~ ��'��굤�}H��q k�`?E���B�W�`D�V�W
r�I����O�!�
�:��ĉt�ՓK��M�wǕ``���B��t�C�=��++�Q�(�SCt��H�&�g9rl	�c'�Ovx1B�F!8J(d;Gj���(���W�O0l���4p�",���>����C�\7uG�C�H��*�=�pb�)m�� Iw����O����hN�lT11�'d��@��'����5��_R���,J�G���ɾ]����努Ϫ������'�ȿ^\�������i����ç����B��f�xEk��'�b� �.���X�'��|}N��-OJ�*S�QO}��U*6�	Ny��9�V&/���B�RLBՁ�"	}ֹ��E�[x����倚�*T!��-}if��6 ��V�DZ��Z�1OLr� ���N�������O�<	���
W�P�B�$��<��� �Tt�P�(�ӹ��\��ھ>� ��L�6R����K
�Ż���1M�phoZv��,�0O,T�ţOb��,	R�
LP8Z��'�Ҽ� i���e��	� �f0`����|9Nߖh��j�/ p8Tm8,O^��&ޖ �j��&�=K����+C����b$,cxސ���H{Ib�B���P��*F�8k���ƇL�Hx�'xJ��so��x�y3W�Z&	3j%Ә'�>0i '5w��m�`C�0tR�³�}�c?�BE �G�B}y�Fсn��q)>D�PW��	>�!N�f�`܋�E
�r���!�����K<j[��<>�I�x�ȟ5�4���H�O���3��\�0?QN�(@��ؑ��+��+'p,�T(�BL&L�b ��1aw��9��C,ay�MR3a�jp�ՆG7Ķe`eI:ՈO�]R��[H���8�X��&c��ۥd�ʤ���~�}�B�#4��J��,4�����=����f ڌH�Ȉ��d����(h�ը��iP��hsg##x��G���ɛ{!���/�X�L9`�X��y <>�M�EL�_�DPqϨ����L�������p<�"!�7b��T� ��:�����z��d�Ige"�S2�\��M܊�� ��X�$5Q�l������ēT�i��%i��Q�@L "�����$�b�O���-C�$�Ei:�i�qz���Ozj������-	U#6D�I��!.��c��#^���sd�d,p!�X�T����@-f|�0�(�,&���4��'��z��{M6e��e��<)r �(4���C�c>.2���VH�e�<�M��[< k��?p��I�l�Z�n�*�kv��%o/�"~b��3�$r��κW_�dg��Z�<I�J؝q�v���I�@4�y�EěA���Ig�Wj���	�(�剁2�F��Q�=� �aL���B�ɜ/�n%	�`R.e 0J����V���֐>�ZF�O�0�`)՜��O�z�$�*�<���b�:n2(�P�'�&�X�@<\n��'� ��O[(7��I���^�#���j�����I��T�@l^5!���Ţ�/L��r� !މ @��c��1��-��S,�F�2%.�6Fq�����H�.B�s�l��SS��Qh�F�W����h>ԛF��6�v�h�JV�O���I�Gv%L�q�c�űt�ZC��6lA�y�pؔGG����#cb�D�F�%�Eq��oDR��韨#>yb/�.l�=2��ز�y��I(<�Gb��9U��P.�u�6��6����K�Pz��ڗR���1ϖjA�����+3�xB�=^j�5ac�XR~���),�L��MU�u-�hF�y�I�^W�(���iB<y KV��)ԔP��&��a�4�<*��h���n7����4�y���Q�`�q���7\�&����K6M�HT˝�q��'�Yf���^�hT�UA�2B���!�'W�=���/2	B�3pL�d������ܲ_e�2��'��q���6\���m�VhTYzϓ^���M$�N�T�)Kd䘆x��p{�)K�=Z!�d��.j�i��E��&bȜ�W��]!��x�.�:�FP<M�8��gM��!򄊧WV�l�V��#W
��KP&�:GqO�-8����0<�v�S�V���c�TQ�P��&�g<�Vc�)��[F�U�V\!���:D ��RX0��?QAN�z���(k�~��iM�'2|���� ��'>� ���C
�ʀCV����p1
"O����]��رQ�J�J�܄[�_�LB�FH(4�:-S3�>E�4��P��3�;O���ޱ�y��M�!�4E@2/�:]ݢF`@����'v����# �ϸ'�T��C+�s(숢ױxPT���=�ZݒA�9%�~�� ��s�a+���5,�k��7�OZP�ek[87M:���(��Z��)��	-o����G#F�O�I���Y�#,��(���.vx�Q�'t�pgT���q�mF�q* �9(O~<b��@�ʹH��|�a��9=��Y�B�>��H��L�z�<a �"'V"���lɶM�65�d�]5��m�NuR6)V:��g�s��lAկ�sw�	UcQ�k�8���s��xq@�]��<	��I�9��رv^�!����o�\���c�2I��@�����I�rD�ݦ�'�A`�G�%tt�y֏SN�U��'�nXqk�S˜Y����E�B� �'f����.I�A°�P4C�Vi"���'T�u��[�����7�D�I�'�U�����(���S1�rh[�'{`��+�O~�d�ůY z�`��'=����ٵq6�h@����u���;�'�tT�����[��`���^�l� Ay�'VF�k'�بH��,�$GI*�����'z��B��6���f�7P�4��'F\,�� � �������K�'�*IB��H"c`�xB�
Ft�����'pH�k�aS�r�K�����'��Xg��%FR\+$�8:�$��']l�@Ǆ�sZ0㴭�G�~���'^�x�F�6i�p��cŋ�J����'��H#�"ΫH����cB
䨻�'�(}��t�:m"���>-<t4x�'�ưQ�O*+����������'�$�r��NO�X��P& ?0B�'�� �@��,��� `�Z��t�@�'td�e�Q�e�dq"7❴�K�'� �i�n�0��)2Wǅ�#�k�'�v �� /�̸g�I�{^v��
�'qX��BH+>�ᒓl��B�&��	�'c���%!�3H@�K��l
�'?6�cڅ`霠�Ҫ�;4���@�'���:��:#�U�֏Z<}>0��'���xu��)!>��gH�kmra;�'��B�0gU ���ƪ2:��#�'��[��ߗ��q[@�ۥ=)�y��'�h*.�=Q��<����;s��T�<��Fo�����c�9w�l��J�<Y��\��	�"(��Y��i�D�<!�~T�䙓���IB�<����6?b�p�V���(Y�-�mk�<9B_	���)�K��*���C�<��'ܹo�¬��*�:90X+��z�<QD$U�gpN0�f��R�i� � u�<5�ی}%��p�&�2A6]hc��u�<qA�
�D��̚�� ("�L�ǮJi�<�V^�b�
�&��Z�ֽ8���k�<A��ϝ ��P#V�L>o&	�qn�a�<a�ށ{BX�p'�3s��M�%�Cj�<!�l5lې��-��q����mQa�<����]�p�Q��<� i����^�<q�'TK��\p���9)��I�	Q�<�GN'_�-���ߝ.�q�ĨKH�<I��M'{��;�,VŊ���Lx�<�w˒�hC<�� �]*Jv8�A��NL�<� �0��E��Ly�,k�<�q"O���a��rȂm�dEj�	'"O���RkQ�(Y�q���Y�K��q)B"O��;۳8����F�_�
&"O��Z�냴N3�M���M��0@"O�p�e�mcB�Z  @}}zUz�"O��gd�.XFD�Bφ!VDE0��	�E��3�
Y���$K+�N�	!|F�9���\�z��@G�"��B�ɛ:��Y�#�S^��EA��I�
�\B�	 ��]��L2����g��[�rB�I�Ą"	C!<�x��
â@�C䉞&�D��
ؓ�R	���_�4�B䉙S}(� �hK{A�
(Q�C�	�t��t��OҷŲ4٠i��2C�ɣIT,ȧ�W���X��瞓k4C��+A��H�O�+�ث�X���B��2M�څJ�8!��H�(JtB��[�A���!�,d7�ԧ)��B�ɛ�u����I^�R SYFB�I�S�jP+6(C�TP��R%E�B�I�~�l@�ug�j�x���BK.�C�	%H�@�j��F�/@�hQ�^=i�C�ɳm�Y�$� 5�Zm8A��|�LC䉧!D0t�J�ns"�+0[�9Z�����l�,�`�'m�lB��K�aG�A�J��`(�O�$0�JՒs�1O>�����,g��iQ�i��4�
"b�O,�z�)ۖE������~*�n�7w�6�(�AX�}�[���B��}{�NC
"���'����	T!_+p�8F��9?S���@�HB��"Wc��Ɇ2I�H
�'C� ����$��a��C��nh8�/PJy��>�L����O�֤xp��	R�������ozs�O6�c3/�S��"N�"|��A��cg^�pEc�֛}�v�	�;*���������u�rk��s(��5���E��X
��
��y�@Ӯ2�j�H�j�B6434e\�y�,z��4Ӓd�?�-�)�#�y�)B�s������8$g+\�l�N���p��q1ϣ�hYX��.F���l�v���k��t�n�!@���<��ȓ$O,Т��ֺ7��'�O!+8����H�S��ޖ �r��S!ۑw}Ɓ�ȓiȽI����AK�]cJF8/�L���D.Lx��Ò9*�\��^�����PT�s #��@�>Y��,��4i��A�=�r�Gaֲ�C6 DI�VI�ȓ!
�ͪWΑ'�,:�DΛa���n%ر�g`\�*E��0��.��ȓ)�����Ւ�x�i�om^��ȓ|hqQ�DԢ�1�.�<����ȓ]>$ �РT��) �r�	�ȓ>sL1�gϘ���gzL��+-su�Q�dR�%��X7Y�ȓS����Ȅ8,^���ݏx��I�ȓ'i,���i�5*X8���M�+�D���$�(���P�A�@�3T�P�{X�|�ȓ��ѩ�F�r=���F��4���F0�pZ�MM/�dy�tј/�ąȓ���u�M�#l5+����,��t�^x"��/p	�q�vn3��|��o��9 �Û� ����O*"h�ȓ!0<�Gȍ�vMp�xv�¶#x�Յ�u�t!�VON��B�C�h|`q��BU+
)%�+dǚ+5E
H��Tq�\��%
21t5�r"�$ԸH�ȓG�������&0�����Y�F%�ȓzJR7���Pϊ��UO!���S�? ��(5�ɡY&���� $]�@8�"O֥�"��%�8�������j�"O��P�c�4tS)��~x"-H�"O�h��#&�����P�Vόm�!"O͚���~
ph`�?��Q3"O�3g�&���g�ծw�T)[�"O����n�`�Zm3��^�~n�
"O���dHV�Ke�3�/i���)G"On #�/�)Md�4���Z�L���"Ot	R�㏣[p���HL�s���e"O����"� \4�Iu��2H|�l�R"O�	2GZe|���U��Ul����"O�,�Eɝ
��d�Fؙ]a���"O=���A'A�|��%H���@iw"O��i1�7˞#ǋ]�y@��P"OhD��Hخ#���	Ak��(��2�"O���.9�N$�t��&���rW"O��B�.
y���^�ZH��"O*qHv�!J��ezÌV�T4:a"O<P$��T���A������"OX�$�خJ���CH��C��X��"O������%�'F�r�䅻5"OPe7Ǌ�R������*�*!)""O� ���P*d)�t
�����	y"OԤ��FT!�(��;]�"O )M�;rT`9�m�(%H�j "O��x�ͧ�ʴ�%l��'�=�p"O"u�cD�� ��� ���4k ��w"OVLq!�	1��	+g@��A���AP"O���s�\�i� U
�%��Gh1�"O�����V��L҅#H�a{�T�v"Oze��V������"HA�8�E"Oni��M��t�M�E.��7�|��"O����W��9�ӯ4^��!;@"O�́w�	�F��pٔO�����0"O����F�h�RvN�(����1"O��C��FC��񦟛i}°�v"O�-�&�P	qM|��%���%�����"O���'j�@��!��^1a��%K�"O�������#�� �"�K�J\Cp"O$!
F�H(q��@�T�=x��)r"O���pjHcQ|`Hq��̄��t"O(�iP�ty ���l
L#>�Q�"O� �@�����kJ:� ��G"O�	�ƭ։~t����	Оd��I0d"O~�Z%��K��M��H�*7�P��"O��b�KǏn?�иէN���ቔ"O0�K��/sX<I��J�F�T���"O�9BC�9��(�Ri
w�9PP"O�����ܲ<т�n�Hq�|� "O��c�H�1�hsmL�mQJ�Qq"O�{`B�0P��A��*"G�� Q"OJ�HAD�
��z@�T-���"O���^%��	�FE0�l!Z�"O�:�ή&�Y1Del^�@�"O��iS�KFk��0 %G��P�6"O8�+�K�,Eh���醎;Dl��7"O�Q�W�� ��[���"l;*�Q�"O� #U�ٌ]z,aCO� ��A)�"O@H5k��OX06� x�	#"O�3�m��4ѡc�<N��D"O�|�F�i�U�!!�(#��U	r"O���	ֵLН`a�wu����"O��+���� 9����E�>�d�IW"O� ^P�W��?h呤e�a��R�"O�}�f�TN�Őab�F����"O�Ceז�� Pdɹ�M�0"O��Q ���+�\����^�0�<�R�'��a��*�p8���,�n8@8��'%��BՂ[����C!#Z�c9�$��'U((X�NP3e�� #�  Eƞ��'����b)áS�v�8��O�:m��a
�'�R1��� �&��ⷅ�0����'��xǡ��0�>i�"�Ƌ}��(�'z�X�O�i�$X���#ng�]�
�'�Ńr.��hA����˝14m�ܘ
�'}�M�cJ�Ԑ��B��&�f�
�'Q���G9qTZL��kR(.F�8	�'����`!X�[S�yC�f°�>@�'���Z���@z2<y�〭(V��	�'�j��5��8<t�(q�J!/�Nea�'�>d�qd�x��$iwKЯ#� $C�'���dk�K��L��i�)H)�$��'� �� ���z4:��;B�Mx
�'A|���B�X�Y�ĉ��
�'���x�뉖���9�!�� )2���'���r�y��)J!n��rl؉k	�'T�|+�d�+%
a�	ӡco��)�'��[��R�u��l����X���C�'|"��a�,ۊp�)�;Ua��K
�'w�\H���-:�" �A��٢	�'�))� 7�T���$������'�ԙ�t�ÿ9��HS�C����'�2�b�-�;h*�K�w
����'VFYC%̵9P4Be��v�JA!�'���ň�!�"M9��˘q)�@��'�T�2 KW@<$(�c?|��T��'3r�Y e�"$�^ԉwsD����'rx����=�������j8����'L��؅��?N*N�"56F���'ބ��� Z�|�w)�$'���3�'C�L�խÅ[��(���N#d��'d>|���_�|�Ե�S`V�G��)��'3�%!A��xd��#(��F`��'{�� )�Pz��"�A�9Jz�z�'�����9���	H|����'`�z�F��C|��T�vޞ�@�'�>�1���+V�A�&DT�u��	�'O�4��	�*	򸘨���oz��
�'h�p�
܏o�
�A�-;5)\ 
�'� ���W��fe�7B�:1|ؔ9	�'f�B��#�z窘5-� PA�'��ٹ��E�Y� ��� �<�x�@�'y���'##F���e��/2��E��'��� 6��e8��#V�Ёt��z	�'��1����C �)lk}q
�'���& ��=���䨎�4�}��'��)����:Q���tH	�,�zK�'�H�avmӽr<D%sb%�b��'�
u8v��e�f�8���*F{b��'O"��a�p�� ���8j�a	�'�0 ���\*(O�t2�e��b�lyh�'����Ʋ,�X��F!R`dJ�'L�L���Z7���w���Qm*���'r
�	g��j�,�Qd�7�|���'��c(hF��ңPn&��
�'ϰ�x���	0��;B%���� 	�'�|� 	R�2�4��nS~[���� ����"�����'����@"O�= p�UN�̬;0� ���<K�"OͺD��b�r��`�+�8���"O�ٳd�J<	����P>/� �{F"OB��QJ	9c���5&�D���Je"O|e�� Ac�>�,�%H�P�G"Of���C�L&� ��Q�%��Y!�"Om�4C_�V��`�o�4P�f�"O\48d�,*N�����h	B"O�8S�שt�a�h���D"O��CGW�� �4
],9L�j"O��q�;L�0��)��iT05��"O̕J�b�n_r��ԧX3@|�S!"O�尢���N]���ˬV�^8��"O�9�� �?�<�B�IV�B�"Otp���j�icbJ_��Pjp"O��(�f(g��p艽'ԁ�"ObY�aQ*��)Gg%>��T"O��"� )�|!c�ĶT���2"Oa%->����wm�.`Rp���"Ol����^L bg��L`^��"OdTQ`��*�ٛ���  Q��G"O  W�N*~Y���j�ZicS"O4�1AkW�| i�W	��LW��˥"O���F�0x��ǆ,~f�MX"O\�6��:|8 �"�j�svBKJ�<A$�ۚA������D�,X(�l�<ib"F?. M�T㒽R�Jy���[e�<����2t�� R�F�l��u�'-ZF�<iу\0gh]��/��Sm@���'P@�<�դ5
DpI�i�'b��щ@a�<Y�J>,���P��.F����Z�<���0k�i�tC)`�Aa�i�Z�<� ��c�n�x$F�(#BP���
U�<a$�	��&aD�o����0�R�<Qt�в��J���ބLC�S�<)&g  (��   f   Ĵ���	��Z��D��"��8�d�@}"�ײK*<ac�ʄ��I&`�r@x��`�\�mڋ3�ޙ� *Z�d<�$!��Y.A>d���41��Ky���5<�L���/�&�
��S�2&~X���04��#<�fm�>mcc*��v&���Gf<ǧ����d�6����*9��	)䚈�żi|����y`��o���p��0t����Di��2������X-��!p��4!S�M?l�:����kA>�� B��)�nQ�qo�H�j�����H~2d��0���p�d�݉z^�ٯ�/.k,S��H1�E��d\���͑e0�ėFR�$��_�<}�	/2��i��dҡ�B+_(3&DX ̌!��E�Q�"<�"j)�W(a M�$��0�J�B�5bc�I�F��� W� ��C��,��	*�Q8n[����%(}�#�\�'}t8�=�%�*6��4q�e��S�x���aɦ�X5�I�T�(���4���C�T��h�L���Jb���S���əZ�t��Nˤ`ql		k��3�ʓR�|"<�P�-���7�n�4⌇Q&�1��f��c��{ቄ~��p� �'\84�aJ5s���ƀR�&�̛�y2��^�'=�%�����,�|���&�<6��EJ�a���j�ɱS�'���	�qb4�{�eX<3�l��G%"G�حn�8lH7s��1A3	��Û�M˄�i�\Q����	�q�ǌ;�ܑyÅ�B��}���+?14oǦ1zJ�<�G;}� ٮ �����i���D�ˀLX	L����^2�(O$��,�b 
6�"���T� �2���'qP,�@ ��&~�Da�Nъ[]<��4�$E!�Dϣf(��lISRD�@���Ca!�$�60��+@ ����,j�L�5:T!�S]�>`�HMn؍���k!�ą+G�2q��A1^mf����]!��C8#��쨶N12G��蠪_0AE!���+N�=��Q�	Bt���א7�!������h2ާ* %�a��&O�!�$P!,
���t	+�p�H2�ݔo�!��,%~l	�/��(�Z�ȲEQ9rA!�E�iBD�I�/�,(�N!#a�PL-!��N>��Hq�
}0 ��$MHy!�d�2^`�D�˫V;:��w��!��S'���&��I�%r�d�h�!�J0Ap��s�܀|��t*���_~!�D��DX� e��`��a�0�cM!��F2z�"@%ѾG݂�@=[+!��7   >    :IZ@-�nkZ��&C�'ll\�0Oz+��AI��e���X�'iD��  ����A��!�!� �Y   �	  �  ~  7"  +   �pA�������\�'ll\�0BLz+��A	��e�2b������Z���'����7�ςK���[4gO�<���V3N� ���'\j��f"5h<�2"�8v�ؘVF�ZJ]���'N]��R�D[�����&�h�(&V�?������?����'�Z`�^��R1������,��'��@�c������ю��횎{2n���D�	:DXL��R�>[��r�z��Az���'T�7�� Ș'�N5�K~�WŊ�~�� �]�<�2Ah�<i�,S�ؤz5��r�hP��
CH����?��I� c�4HPF3P|hx��W{�<1���}SrJ��ͲH���f�F��|O���7�Z:���(&_���a(�0i��$� i{���<1�l��?�	"A�]����v�Y�d�J�6%�E�ZΪ���/�3���*.���1H>���I�Ut<!�$I�S�}A
�]��a@ə�l"1OZ�=�|�qG�E~�V/��Md��ic��]�<��-N���d�E�4�^�g
�(�HO�'71�O�JCh
6�� �bc�G����'�����6�I��"|ڧ!�gBrhȁ@
��F���6]t�y�@NU��8s�G~�b e*ΤC�L��#D����U
s��LöNK
;��D�E"��<��œih�l��(R����Sf�<�d,W2^��5[MΘr .���������O:�Ez2�0�$�9j6�b�8nYtm�m��UQ�!D����ݟ��Iџ<tL��Y����I�|ʗ���4�$/�0ϒ�J� d���KS"Ix����DG�t�R��'HܧS�N ��=(�2ԨT���.Qbm��E����J��QʩZӉ�Ɵ��I���	ky��'��O��2`,>0W�]H�4r�{s�',��O�H��N�b8<�tFR�6�X�C���$��d�<Q1��6M�򤛪�p<��C�t{��a �L�0N~uJ�>���[�Bx�OT9�!h���'�$�r�f@�<f��#�����p��If�zd�|rm�"*��@�aɐ�EE��°<�@����	@}�@�fY�Tȥ��>n���j��~z�������O��%bD�J�;_�xۃ$�{wDȊ��$�S����t�~��wg�/w|�	 ,�$�B1��'u�I�!uh+�� b>������B9a�+J�@���%lɾQ���v.&}�U
)d��c�)��M�3_��,��V	�,	��iL<gbO����)��9j0�@�+_����KI(P�pO��9�'�Җ�ԙ�4f��<�)�`�M�`HPx#��ǫ�(OL��d�[�P�!K�V����n!EZ#=�O��8J�2a�N������&Q�pVK*y�@7e�O:���Oԙ0\{_����O����O�E�
�*S����JÇI����F� ����sc�$|����֩A�U�XC,ׇ_�S���I�hX Y3�R,N�9�ӈ&j�U�����]�����M���[�ҘO�<ݛ�,v�}�-�1)u��3�E�h�'i����'�"FU!�O+��'X��'T��m����A�M�	P�N$ s�K�S�4�?)D�NI�h�c[�gV�-JRFW�����I��yB'G5�yrd����ʷE��d�~�aQ�f<2�1��ޟ`;Z��B�O k���8Ǥ˿=!�Of�c�.�C�AO�Q���8i帨A� ]�:*z��r�|<����;���)['L(�	y��V�2���8�� ��ЏZ����W$U'&֘�z��DȟȺ�eP� ��2�l�p�@4EN����k$����P]�@�҄+V�[�Ҹ�=9�Ė��Tu��3��<9�4M�`yX'���o���&[�Zv�A�T�'�B^7ub�숱�'�2(�$ Qx0�3��yR�i�6�RO��N0��sDA�]	 �	˓UdR����L�=���3�E�O�h�Bg8p�^�3`�� 5�`�sU�'������?���iۛ&b]�j�:"#����D�Vբ"���?ъ�OK�'�F���A�fѪY��I�>ȋh��|����'n��O�.�H6��
�ͻ2DИ�?y)O �Ɋt�`�D�O�˧q�b$��4~��m'ؐ��!�c���2�'��lP}�c�]�>f��v��O����+����'y�L��ǝ�D��D��E�"�}%���C��6�H����,F�
�*:��t�q@D�7�%��CL!��ul�0�����F�d�i��Y��$Q1<L��0B�������*;$���Q��ߤ$+u��R��h�Z�'G�)���O���􌙰a�=TB��	!ֱY �Eo�Iן��	�p3�D����x��˟P�	�L�  #�=`��;5��8��e:�"^�y���'}Nu�����A;WkB�i�Gܡ.ı�>	��]X�̠QEO
�1��W�_q�1yË��?��?���?�}���C�ӗWRl�Aɕ3`9�K���;p!�ϐ+r3(]	L����W�W�#$Gv�h;�<��?��������:	 hM�3�J�s0N%�(�x�lT�����	�����ϟ�f��,��d�	�|:ӋQ0S����\[�\�g�q����J6oO����*�
�t��t��	Fo�5^�ތ�5)��q`8�Z�i5�OH�Pj�?1�P(�!�� ���U�EJ��oaӆ l���'���Đ&~� �a�dƘS�rQ�d@�R�{#�d���x�t��1�Ebt2qO�L��6O:ʓR+�`z#IB��?��4h�P]z�/U7b1D�z�F�P��F�'�R��3g�L���'����Q<�!:g��yB�i��B�o�c����f� (�t�������R3� Ё�O6e�֩^�|��2Q�@ ѫG�'
����?�E�i؛�ḛ3>��)��Q�e�C[�SY���?���O��'.\}�P$Sp����
q�J-R�B�<�S�EA��̬���?2�y�P��3�R�0F�',�ɭ	m�6M�<�����1'.p6M׷TȾ����G�Z����׎C]�I�����`%��R5b5)D�;}���*�ӡ΄�̪1nH�~@\�N�d���ҋ$�D�
��m��B�����(X#C�	c�P�$cǔ]�.3��xbi��?���?!���Oj�][5��?es��)@B n�l�0�{�'�ayR�U�NF�D��4ĺ����������'n;P,�?���޿B�ee��7g�I���=O]�ѩ�'	�'�&Q��J9���'��'>����)>"2���n\<^����S�]C���kJ�p�f��$�65 ��-e�v�;�@��8��5p�0
�(��%.Ye��Q�Vf���~&�Z�/�~��Q����(Id��s�D��?q���?��d��?�}�'�FƗ�x�4��s�	�s70y��K��dZC�,6����H~t�e���dR�<	��N�'�n^�l�'Ѽ��0	�kz&�8�hƂ		����'�4���n.��'H��ÎT���Zʔ���R��`_0z݅�k3Rd3
J$D�a�DC:pVA�ȓr� ,Ce�E2����a7~��e��'��D�������'C�mD�AߓCl�'�����e�:L�p��dDa�Ę+��+#��:e��'l`+���S��#fFS�Y�J���fF�b6Vc�<��?�)K�!!��)�<LIS"*X�4�!�IA�p���E�F6\��NI��azr��O���|�Ì�1�T�!D5L8!��¶K��@qcE��h*��; O'n�O$Fzʟ����h.V��ؙ$LD�	�=��C�'�2����(�Ɏ	�����*TXc��t���s�ʛd��b�D��!�O�q��'�y����F[�,�7Gԩj�M��'i���#�><��W
��S��1�y2�)�Ӎ�~���])����b*'��C�I4`�t�C�$Z~�� 1+����Fzr\>�+ǿ.�d�I��e�1���?���� 1O|�!ᓓQ\aYq�V(T����L�P�ҍ�)՜����y�2��B�8���Q��čz�!�č4q�:y��%�C�>Lp0�j����� ���A�����C���6��C��?I�4�x�L�+�4�iʓB���k}2�#�M�'h��D�R]?\�#ζt����'�}k��'���ƚ��NȤ`L��6�d���H�:a̙����f�
6O������4B�T��ȓ��q�U+ɽ-��r!�-h ~):
�'���2�$�8h����A8)���ߓD��'[���ݡMSa����0@$`�ь�)ғC!�*C�'�#�
�������0v|��YO� #�IB3S��b�,;5�.�)���䱐Gͷ{�l$(E��	=G!��m����ߛ{���Bό�p=Y��H8&�vh姃*4�p��J���y��Ȥc��T;T������#���'��"=�Olv������|Ȕ�I�	ȟe�^c&�8�z�,;4󤈩_�$��5eN��!F����"���1O�� ������S�? ��ZVC����� �-��4˜�H`"O4���o�X��C�Ï}U�j��6�Ş2iH-1
�v0���Pj^k�Ņ�2FHHT �H��PC����1b�����|�"���g"y@a�G 	�
uӁ��2�E�k�c���-#§]���9f�̗sJ�H���f���O�c܍��	k�"x�D�E1>�y���34�B�IGV��:�T��>	pAg�<R�#<!ϓt����M�])��ᭅ:#�ȓ|��܂���pű���3^V���:��d�r�'qZ�O�8� K[��!�	�/ܖ�;w�O��&�F831O^,3W�FQ�'��P�#�!��0Xg@A�gGQ��'�5H5O�	^&�����<sϴ="	�'{}���YS�E�o���B O6����:������	����I��'/2�O4��c@�vB���Q4#m�*A�dF�'e\Ѷ��O�EY�N"��4+��+NҸ� �>���3V�B��<��_k�S�jk�@pS�8�����Ça[�C�	6:u���N*�C�FOQ.���9��8��eIw�W�o`��3�m͑mB�	�~8L$y��< ur��!�L'��\����?��c��0�&hX��_0"��|QSJ���HO�3F.�g�i�����&�P�1jUqa�����X�~�rm�<��lɃ~؀�>�O^�a#�&��h�Q��H�!��"O�Uځ���_� b �B�6�3���/�S�'2"�r�A%P&��E�Oml�ȓw�3�Ċ�= �h�W�
�1��`����|����ֱ���	�$ ^q��F�3��LJ�pf>c��J��6§Wy$���g0<�����=��%	$C�~L���	�E��1�uC�;}����I��t^B��	s+�(H�I$��MVC����"<����Y0��6�p��6{�>Մ�P����+L6.E)��2y0�)�I0���|�'Q�O�!(t
ފ: �!e���4x���ON�@�ӦW$1OZ����8��';�=�OC�T���:�j��d ����'��scjA�uB��[�&ƲK��a�'�E�G/ܦb0=hT��>bnA��O��@s�D��XD`7g: f�Y��'�z�O�X:�i�y��D��e\�r��;a�	S�'�F-����O�PCr�T���	`�[���y�>��!)9@�<����E�9R��p�H�0A:d�Έ 6C�ɲ2� �r��/4d	���ˋA}���'�I�l*�ۡ���fh�L��b�+��C�I�d}��Y'��&h�|h؇�^�E:�(���?��b�1��k�-	45:L�����HO�����g̓
���}���f'��3�L�AF	}(,�<a���!}r �>�Oiq��]�K���p��-DY>��"OR�8�K2v(�H�"Y�p�Z����6�S�'6�Tb���]��A u��;J ���fg�XH�$�m����9|�r@H��D�|�'��ʄ<��P�pkI��i��1+�g�*wH�b�H2p((�'H����6IG:i�(!�$JƁ::��qa�P�m|���	�P���K�;9B\��f��	FS�B䉪6�@�bd�6k�`̺��%� #<�ϓ{;������><�Bު:P@�ȓq�x�8`��#,��Ԋ%�[sr,�	�����s�'�`�O���C�z܁����v5L��S�O��2��*Z�1O�9��44ƒOZ�1�A��ZPZ�J��S	��{7"O:M3�
m���	�ju�"O���[���`1�Z
d�m�D�!4�$�W�؄y�x2�Ö/�� ���5|O��$���&<fl�4�ף(��}	4�	P�'�F}x��O���@ ��f��IZ�j�B��>���ۋ\���<ApT��:n�pX����Zy.9IR 8"~�C�)� ��M�,���q&�?f^�r��'��OV��i�&�L�7�ڿQ�B�"O�����%�B��j�.[oV����]J����49rUF�\��xP�6o\�EGzbHZ#sF�b�|�g��:�2`̍NC�M�1O�.n��ܳp@,�Ɏ.^�ݣd��|��4,���2t�׍`���AG)�y2��o5<�P �C8
`Q����'Eўb>�P�C*d�1�*�U��$��(D���Ul	�oJ*4�!��,@�3.RY�'���'�LY�fGL09|(��`h��z���(�:�h4��W�>�H�8�x2�厈6
X�)��+��5l/�O~}�rC�2Iqz<�0�
7x�h�	�'�� '��8e,>0��$�@�R-���5<O�ڤ �"cbn��7��6CX�y�"O±:3�܈f�d��@:b
 ۧ�'���@����K>M�;fIk��B.��ZE�T?�#�{�č�<#�'h��$���nĲ�xX�G\�In�jUA5D�P����.�Fܣ�l�iz��!
5D�dzF��m��аTbd�ڕ4`�yh<����)�,�@��'7|�q{��_��xxO>!���9��ac3ǚ N���QK[�b?����䔤�?)�l�[�
�B�N]B�Z��"}����@a�R%7�ODr���W3ڹ�bAX�I���'��i��K;m����`��;+�i���'�,��$^*3�$*���#;����'�,h�jE,ݛPH�eR�1��d0�S��01C~e��ĝ-�J�Aݓ�ў����/��'0�����!2�AD�?4b�9 %��	rT�y"�)>r���}&����K�����{9�
B)Xr(�B�I�LŦ�Rc��8gk��X�ךS�hc��F{��4��J��5�R�T���mQ C���yg P�:,��J�^�Rt�&V�� �O�X�\��lY}E���Ȕ9༜�Q��Oh(��Q~�*L��G�T���z��4��`k~$b�%;K��$�3
�<��?I ���y�Ϝ:�j娐W�<Q� %�ISS��$KnY�Q�EO�'��y�O7����T�z��(H^���'Ԏ�Q�,�gr��D�1d�"���eI���HO��$��B� 9C��2cI�*�b���D�����T�4�b��]�tm�O4���-ř
��0{1 �=ƺHb"O�-��k��{�q�.��s""O��f��m��J7N���a��>4�P����ln��W��M�l��w�:|O��$�Th���<t�ιj�:��}���%����HOb�H#���Dʗ�88�&q��,�]RR�:7J#��m���:�y"�I���l7n���!���#w/Y�qQ2	��dBI�P�ςF��|c�ͮr���	C�W�8�:���V*�Y+F�4���R|zq�W��9q���S�B$GG��?���)��N(:;���2N��7���30�hO��[�eq�8@���&J�*�``Bv}����	6�l�<��	)���>�ON�C��� fA��e�N�*4x�9"O:���ϐK�
����J�,{��;�u���O�P�۔'��T�5M-����'}4<��ԣy�6��FW/d<t���In�4'&�	0"��� Oջ.�,D��
��:���.s�@�<!$�(�矜yq�K�&����V�/b�	EBι����ɘ��#�-� ?���S��Z"L\�B�Ʉ
X(a#2�X-ʴC�'<�"<�ϓtX��o���4u7cƩ2sJ}�ȓHvAzEj��SC�Lj��  �J��	���dBs�'�1O�P�B��i=b�'	4���Rw�O�)�$�A�1OX(�;8��$�� �NM7���r�Q�4�B&b4D�`�Z����P$*�H�%�3D�� 4�B�dD�|���$�B"���H34�Ѓ���Dd�;E��8L��$/8|O`&��sA�H34����`��P���:�I|��u����?Ʉ�Ý(F@�����<%�B�3n�I�mc�`� G9����x�H�´/�
k,��9 
!�$-\�X�Ip/�0kL��d
m�az��DI�RK!��L_� ���6:P!�W�ȅ���` ~h��.�;:��OڄFzʟ�d�կ9� ̈��Q6ЭZ��3��P��d�����DǜP�2��f�L<!u�1OL=)3���䓄}4�.I&UN	�*�+}.!�d� MO��91-��&qY7���|�1O&�=�|j0k[,CE��!Nލd� 6�[`�<�@ި�䀣R ��6� �9+>�HO��'0��O���a��U�Y��#�:�h:�!�o����O���J%<�B}m�՟��ٟ�'��i���?,X1�P�ՅI��#�C�;ӌ���O���3(���4]�L?O�̚$U -� ��	QL4!RC�jaȁ�X��!�Ċ����8lY�NM� Ð�KITI�p�'-�I���4�2"=�U
ŕU=6�'��r2��v	�O�<y��<�x�wmҼL,���BP'(��Ɉ��OZ�d�>�
1L2��GB�s)p���͜&Ъ��gaӖu"��O���<�ցH&�?Q�O�&i� �(,t�#����j]�ŠGB��;}� �1FS� ff!�5�S�NKh"?iQ�D`웓+_�T�H({��U�o@�Y8���
�V��Kʫp)�Q���	�l�dߐV`�ٓ��4b��i����O�d'ړ��'H��"L��v�j<�5m�I
X��ɳ��r����I�t� �W
p'0�=�v$8�?A,O�@r��Q���iB}0�B���b�h��Q�HK ��OT�:F������dΊ5M��`�m�*1�ʈ���	�D��D���Zy@�.G�,t���	��Ȱ��T��X`�q�O&f;b���g�a����t�x|
��'��?Q�OR��wC��JP9u�%7lH�u��/lO�T�i_E��"�������S���I�(��x`�∧.���#�!в1�ङ�*�O.�@�咓f�G��Q�����	^����;@� �г��B&�C�)^�x�x p�'["eX v<���O�)d��t�Pc�O��!N�8�x��"�4l+n��b@��0�l�qwQ��(*�H��"��/����{�Ob�92�E��4���AtlK(V|��L<q���ޟ0�	u�O��G�h���y$#ނH{����)�y"@�aSjԢ�O΢?��
�	�)���L�'eJ(��?�֪�P�ع�+�H�s%�C�~/8
NS"���'J�9�֢s��)�O��D�>aB�	 lԬ�T�U�pMb��)vJR��놊}ۖ�?L��%cV� ��3��
�$81Cp	ւx� Z㨕-J���:B�Z�4�������}ۧ��x���+Bj�IA�$�F%���J�T���� ?q�ݟ�M�'���s�ǜ8��|ja�!��5K�'�0��0��k�����t �	��yB�+�O�$%�O6�Ӡy{wLE�]�ڝ�q�S�X)6�%1���n���I��'�ڜ�u�'i�X.��y�G���rsn��X=o��A�n+��C%!�I؞ ���u���cb,8� �k���>'��L*�iM�(ky��J���c��ʍC�/p�xE)ã������u�'ѱO�Y�n��ݢ��V�΅y��a�'�O�]#B��r�N��Q�f����$܌���9�i���b��~�s�$U�<�t�K���.:�Zv��ۦ��'q��L~$aʱ8��y�N�'V���\4�B��=LafM{D@�NB)����;����9�	2ԍs�a�O�x��%Y*AunB�ɑMw=��ԸP@��vŗ?F6������?�O�b������]� ��iȲ��y�'g��:$D'��2+g�|�h�i5Ǆ4��� �eZzb����%�q��'�<h�� �%4�f����ӷFH@%R�'�8QG�͔IC\E�EF
�0��y�)�ӣE���g��"7��Z5Flb�B�� (Δ�:�/�7t��A�OT.�DzbW>E�B��)ID��
��H�(cd\��y��'/�p� ��   k   Ĵ���	��Z��D	J<��8�d�@}"�ײK*<ac�ʄ��I&`�r@x�`�*�m�5J��D�kW����`��X�����4\����z��u��I�v�"�]�AH ��`G�*yPTAg�#�U�#<���b���#c�kZ�z��\W�0��P_��0!�˹p"Z��k!?�J��s�7l}2�G�Z�X���	}����W�E%l�L�h�녌,J���O�<�eB#����Ҥ�O��S m��3�Ň?+��ӵȌ& ��l�V�^�l|��O�W��=���Ο����kݼ{��IhYc�^TQ�U���1����0c�g?�mߕD~�h��L@~��voڊ��d�d�֤�p$�*a�\R��У\��R��O�P�����0��pg`��sZ�������GxRXI�'����'�A�Ca��A�BH��őI�H�N�x����omqOd`Z���\�� c��#�^�Ƽi�R�Exr��u�'�ά��Þ�t?ځ���& pM�`dڠ��'�8�Fxr��x~b�9m�l�;�D@�r�L��f�ҳ��ד�O ����M"��R�3px`�����'�|Fxr�Da�'��a�I�p���-L�b�C��k�Lb�䠳ታ��'�����(��I�F�a��!��'9�Fx�/Gc��~�F�nl3��95hh�CB�| �F��F��ɀVqz}ps v���BӈX�F ̠os��N�	�b|:�~ P�ȍ�?���z�2�"@�$ʓ}4��'^MjWj�����[��O7*Wd���ȵ(��)����O��CV�,��W[����"O� ���  �&��"O���eҒ2KD�!��~��S"O�}��`��]c���M&&ظb"O� r2�%`k����ω+o�@��|��)�.��)e� *:~p
6�
�r�B�ɂI�l����J��Z���	JZRB䉥(@$qI4N��w�l�%G�GB�I�D-f�hT�I�H~-[���7<��C�I�1Y&���N�%Pt�ABrb���B�	�+|H��	_2BE����Fw]�B�	�����e\ӊqe�E%DlB䉨'{��3ʖ<Q�l�bS��*1g�C�ɠz[ҭ�i[0K��@��i��x1@B��0lDC0j.a����W�7Y�B䉒)b~��'� Ni#6�1,�*�����'Z�R�f� :���ɔFT:FC�	�z.5ku�@�;���҈�4:86C�	�9�T,�   >    :IZ@-�nkZ��&C�'ll\�0Oz+��AI��e���X�'iD��  ��J�p9�l5D�0P����   �	  �  `  "  �*   �pA�������\�'ll\�0BLz+�X @��e�2b� ��/?~��'������m��.#���2c���JW~x���B�n�HJ�H�#?�J�+MT<@K��xx�P[���(�P��K�*2�艸6�ױ=�0�$�O��O8�d�O�b���v��7_*�s��I�B麽�W+|O*�%� �s�â >(B�"ˤD�
��$�5�0�M�	S�y���r�O_�Ճ��j�8��f�J
@ <QJ������c��C��"����d��C�Yڀ�4'[�n�!�d�>8i�郑�K�I�>0�1G�d�azb�DП�x�"�I�j��}Q�Ȏ��!򄛁_D�S`�<���AA ';�O�EzʟV��,$�$�l�+#�V�Ka�'ړ*���0��䝞W��DK�1�V������,1Z0�ł��s�1O�����R����`p��(�e����G8dK4)�ȓ�)b���b�^�r�N�>����<y�����"Rz YbC^V�t��GT�V�!�$K�`B�ڢ/N&LdT)�1$�"=9,�(�?���^��1u+�Rr�#K���p�p����'+ҥ!��;F�|%�pER�3�z��G�7ζ�r�עM�"a����
5/
x[l	��M��y
̝ZdB�+���$g��=[�ι�O��dO�F�q@�K��ƍ
���]!�B�o�ʭq I�a�Px�Bʆ<]��&�>�U�	+��V� qP$C�sd�R�����a�(�+� �C��'t��'��<v=���'��R�'5h!9vnU�	y�e�O�(3��aO�e�1��d�V$ۣ=����`.I5!�DǘP�������Z�p��J!ظ���'�R�'��R�4��W� G�p8��JY�\(�cJ2�>���Ɏ��vR�Z�mC�'�<�0E_���i�=�U`_�?�.O�] ��UA���4�>E�X1�v]�#"ՙc��TW�>1��E�3גɦO���fC%��'?�8�p���3V�$ZQ��@+Zm�剕]Sz `��|ү�V�a�vl�8L.u�"g˾�<Ʉ�֟��IZ}rB�Z�J吂�$7���ps�ǋ�~b�'
B���z��̆�%�4��qoʉk�1q��J{���)ˉ	bT���X!���`܌%yąyc�O��U�X]!W� gj�|�����u��Q�.	,��D(
�BCK��C/a�\Q�e]Oܧ��By��^=qɐ�1"���]f�0'�h:@�6�S�!�� ��è;0�b��W�Q�N�&�lx�$�Ob�d?��)�~���!�N�L�0�@�`Q�Q���剳M ��-�u�"a���_]9��Ez�؟��x����
8�
 }Pl���T�Z�"��Z���IƟL���"S�	�	ڟ�����ܡ�käQ���E�$�@�*��
N��DK�bD����������$Q�d�'{� Db�2���c���Iq��,)�t q�X00�
�� $�>���M 601�����ۼ#C��$���n�XO���N2.6��O��d� Sc�4����O����OP7B1�,d��!RCC�yS"#ݟ S  E�)�8��'*~��"��q�8)��Ɉ3q�8��0_��W�E���Q>,��	�i^��x�DF�\U�`3���%�����MDdJB��F!\d� S��B���'��0�j�}:���CG	-��Lpƌ��x����s�����#Yܔ�8��ƞF���'���r5k�]LV���U~I��*�0�?a��'L��ы	����3�O�#Cl"�1
�Ra�'�����?dCP	0�^�m��{�pf�|�LR�G
H��'��F�Z)����C�� k'�H*p`������O��S���26l�$�O���0�ޛB0��9O07mR�z�p�3�jIw�p `�3Kay"&/y
`���W����I"!>�8q ګ.@�|b7@Y,*�����@4Hn�'�7�h�\%��F�9�s0�� �`p�UCyb�'W�O��(�DR�L4)��c��`Ɉ��փF �O�]Fz���0�"cŧA���;.Ā��I�3"��&�'��l{�����������2|�6!�2*�Z���	*^���hݤ Ix���O���v�Gxf
5h�EJ��F�韠�dDݚv�4	��mG�)2�EA�B��Р��W��7�����Q�/���B�Ʀ�(��h��CڭD��		��!08L�:��xbh
�?���h�7��4<�䬟.F��A��\�Z|��@�H)�'�ָv\ =�тS߮X��?�Y"-.�	�cH��1��=�!�B�b�4�9�e)�?���?i#� k��xZ���?����?�F1�  $���
eP$*�I�+jd��R2YV��'˓EH�}�fGB4r|��s��X�=¬�>)��]X�bO�����\�F�)�1C�!�?Q��?�pğ��?�}����Ȝn�����ŷ%��@iB��q�!��KV�.�h��,C���i�dO?Q>R�e�0ɓ� ��?=����䝒�l��q��)I�0t3�חSX����A���!�O����OF���H�JY����O�S|�6�[c��#H�7cG�U1�4�E흦1�!�f:�O����#������=eI��b �[�KK����?N�a|��^6�n����٨1��1�`�րR m���֣t�2��<q����'j�E��%x�sĊ<Rڔ��(_�'KR�p�<۲��5@�#/|ʝ"�{#N��y"R��a�I�8������ysS�ʭ*�Rٙ1-��Qk.-�1*���?)��{E��x����?əOȂe�S�ҁlʽ�'��;�cX�w�q��W�Z��Y��dB�k��ܺ�dP���sGY�¨r��K&A�L ���2h���O�Dj��Yъ�D��x�c˵�$Y���@[y��'��O�\����;�b���Ðf�1�A�d�K���	�B��G%G o�
j���LI����<��G�;	̓�?9(�5���oӲ��� �ML�����§x��p���ʟ��IV�L�ᦄ# zӧ
�ĉ�)�d�	E9vdk�ș}�i`A�4)�Ox�����A%�x���i�(X�J~0qdj�?*����x����?���?����O2Jlj���0+��,���ڤu���{R�'�ayB� �{7T�A��:9p��[��O������j����?�#��Y@��A�	rHij�.ϡ�mP�'�R�'Y��󬓂fUB�'��'.l)0"+��}P2-8%%Z�D�.�GR�1�~Q�N�C��^0fA3�퉳&㊬0'��_�JL1䬋�M~,u����S��S�~���~&�����ʫo>�5U�D�rN�p��9�?i���?����?�}�'/�f�	��P�&GC;U�L@q�ՕL��B�ɅN-����+�Lu�fD��<�D��<A��i�'E������'�r Д.,<&�zs$�1h����'uT��.$ܘ'������_���z���圯O��z��=+���ȓ(�R���+���I6�'���ȓk��d;��ލu��5a��Z���	�'���D� �^).�1b@ٙv� ߓ`j�'�L��a��oݶ�g����u����"ғq�4�r��'�퀃jY
0���1$	�wu��H���P�V�Pټc�$(6�$�iS�D�L雖��b�Rx���ߨ=!��)gt	 �_M�`x�`�U�az��Ę>{}���K�c��÷��!���uQX4����(ӊ���Ƣ9k�O��Fzʟ.�� ���Z,hG��إ��
V�'���g�'��i�h���1R.�
���.T��`A�5r��c�<#�̵&q��'�V����(sR�Cٰ�'�%i���$\�kd� S�n��y2�)�Ӈ	3X�s��%U��IR	pG,C䉣@�����&J��h8�`�VQD�Dz"^>YʎҢF�\k��Z�针!�T|��g� �?Q�Ze1OQH�����M�Fe�B��0��� b�2-*���|���$ѦL�B����XǴ!�fd]�PQ!��ك;H���,TZb�l@�H�,��ɜ=�0 i��v��<ArD��B�ɭ}(���T@�,��x󣀍qF
�D�B}2B'�p �'"<���Y;[���!��"l��'�R�I�꛲Θ'��]�W�BI�<�'��E�{��W'Y6�--D���	�?r���R��>(���,D���"���֘I�H�u�F%S$��eh<�r��zzh��������X0��]��L�L>9r�J�C���"�	T���!^p�8[��ܣ!΁�?�Cˆ9:�(ɹ�C,_ܴ���Mo��_�. K������O�X�k�ä4��}���K�;ހY�'��5��k�(�G.��0ȼ����'fB��qےn�ҭ���F�'
����'���aюA�]�]JV˗q0���R!�S�d	9B��3l3�D�kD�N9;^#=��f[#u�1O@A��OUC���)<,��N �|�����3�||���L>� �p��		�Hh�w��(s��R�"O�� �
�5��,�c����,p�D#�S�'!�L�󄞱���,ա$��ȓ{an �"!U�^���#x`����Ĵ|
��dG���+�!^�D.мK��5�bO}�b�<��m9�'Y��!�J�T_b���ĊDWڈѴ�G�k'L��	G;l<�����j�V��W�@B�I��4!k+�gb�����	K38"<�	�_��%X�ꗢ){���F%7#�i�ȓTo���5�UV.��L2\�Bt��7��d^z�'8�O� �&�­4s�e�ԍ�X �d���O������1O0��̈́��'R0y�N�"t�u�p����
�'?��J&�~	x @�ȕ2�4�P�'r,�"EM�VW�}�&L��52�U��O�a�J�1�䐑saU�Z��4y��'8d�Ox�1���y��`LΔ[��d�V�'Ƃ�� o�O48P�,֊D~>H����"*9�ؚs�>qd�N�E�0��<�rg�n��

x�c�_q��A{�J��7��C��;�&�T�M�e�* ��f¯.q����7�I0{�U�P)$_Hc���X=�C�	�5'�袦�ֻbf:�k׫	�d���h���?��S(Y (zL�قBS�*�jY�f1�HOz��c��k�^�zQ���XV���Va�,�uL^�U~��<	�����>�O��E�|:���g��,��D"O��bCU{fB` 昦)i|@r0�7�S�'v5,��2����£�[Te�5�ȓ;*p|���\�">%�fȜ�!����ķ|ږ�*i�"�8�暭
����ʯC���1<�Pb�`��%/§�q㥭RL^\���ߚd8���lQ-^A�ل�� ]Zj�SA�شC��TO�=�C�	�$z� �PDŀ6���؄�Ĕf��#<iϓq���r�H�0�� C��	i7���2ǬP	t�H�j�f$��͖��	���$Lk�'I��O�bB��]�<9D��Y�:�y��O�A��a�m?1O�X%o�z��'����c��	S���1��=%�ܚ�'u>U�c��6��͚�5�N�
�'���9���g��=XgN"_)(p��O.��0��$bR��P !�'�O��K���	�f�eG\kT����$�a�'��L@��O,�q�aʤe�E�Ҭ'��[U�>!�D�1N>(�<�ae�j�Aj�0� Z"7z�)bF!A�sȆB�Ɏi7��H�fM�x���� a�z��$=�ɚ���c��V��2��@��*`~B䉏`il���*��o��5I���
GH⟐����?q2l�=@ú�� ��Y)�����HO���A/�_�/z���9Q�h%�Lʁm�|��p�.v�L��<�6�/v�d�>�O�u�Í�<��5
0�s� ���5D�P[2+zk4Ys��Tڒ��M'�|���O���{��I\m=Z�9f���'�L��ơQ /�=��i?-�	��I\�4�1�I�T��Ł��3�ˏ���D�%���<ac�S�On�@�D��)�B�����X�<"�,O�y4<tJ�JJ�ͻ2;Up8�g�L�h�rЅȓk�}��Ҏ)F9{T��	Exb�'yp4�2$��E�LУ��*��' �r�&ߚ�uQ���>�ܘ���k�I�HO�l$��b��L�
�0���� ��ɧ�a��Z�9�c��d�i��&�l`�CJ��,0��.�W�5�j'D�<Jpɒ�lyn0{��Ĥ��qr�/)D�x�"�*fl�A"$@�
(���o�ch<�e�e����tc�:i��[�II����I>�P�ҏd�ZT#V��9e�F��bKD��hO��Fʝ���	�2r`�����".#`$Z��!}��:\Qa�y�B���'@���KEAF=;�~� )񈄅�S�? z�ض'V�u.�q�@F
A����'��O8x�ݫ~|��JC�N�O^��G"O� (�$�g$8�1��$"j赣���Pw���Ɇ�;��3�P>yx�¢���F�DzR
��c�XA�%�����U�@ϒhR�.!T��� 0��:�y���|B�4=k,u�c�0iT��BC/W�yBi�R�,HP����#����'�ўb>I�6b7j�Jl�#�VyTƨ�A-"D���U*��'qF�2���_��[գQ�'�S���'��0"�*S�"�CWJΊ9L�Y[�zW|��2���W>!)�@M�u�z:0댾'.���U%HRK�UH�''�O@�e�j����U;@m�p"O
��匸p��7��f hP�4�yx���7��Z@3��Kl"<K!$'D��+ �4�~���.2����h�O�Y�'U|"=��|R��1�,H	'	 %��=�H�~�h����Ղ�yB�O.U�J>� ϖ�F���BS�0_̄���W�<)�DU�[�P����̺DԂ A^o�<�tfU�-�`
d��_�V����Y���x�@A�5\�,1C|�3�Jg�dP��I�����!�?7��(���&�@�?A���<Y>���Rͼ�c�� NP%B0+΍>��E'��Y\>��<�'c���8�3 O��^���ߏ|��B�I�=��]{�T:]jW������$(�	,D�����5FE�a��KBC�	ciJ��#�RZ��83wN?������?��$3&���cT�3�a����c�'�x��2c6�ɪ �x�i4�h:���k-|�ӆl˶sZb��h�Զf�q��'� �8W� �yTHp��CK�\�(��'��E�0gǧ�j��3�\=4��D�y�)� �N����Hj���Q���B�I,$4�Ԣd�<�֩��K\5yzEz"T>����+T�!k��چl�J��D�?ᰡ�yp1O��G�S�p�8s�&n'��P�l�8}���炞�\]���ėM�(��!� �\is�نQ)!�@<K��m�c��a!<}h�R{����	$T�� 5-��.hZ�OS?D7�C��o�90���U����3-ɚ���q}B&4ғ^�'2�QȒ:	u�rn	�A���'F8M�sG\)�اuwg���tV	İ��s@�U�J�ȓr�J�o7Py�Ȓ���.�������Q���jT��8�j�,E4�
�'s,��]�v��#�(L� ��\�'���� ��Fq��ω��f����-$�t � X�'�z\���)p����Y>i��K<)�	�znb��P��2�	ϐ}}T���i)ޔ+ŬL9(w!�D�G2j,���E�?�j��KO�z\az��Q<-@ !̟�{�J�ض�N�H�!���y1�ի �ՎRx�Y�A�� ��O*iFzʟ�@���~�h�6�MqԠx��9�NО��r��
��ĬڐJ�x�τ�7�be��M�y�1Oٕ��)ɸ��GHe�����4��1�*F c����g�=�A<W���x�H�$y[�Y�<Ɋ���S�##n��AE�d+r-bӮ\�N�!�fڌd������2��N�"=�+�4=�?���OF�U�G$:sp�Q�[ڟl����:��'��lE���/��hQ㎋1�v!�$ꉚ���A���?I5��6&c�͘�&�*r?��K`a�A�<	���5r��P�uͶ 3�W}�'��y�l	���׃�7���Jw���y�N�!3Z�Zr�20���aO��?��Y�����,�%S�L���R�K�r�����"DՌ�I�k�1c+执�u����sD�(�Gm<��E#&�͸!�F���y�I�!Z�`�2t�H$Q����S�? ݓ�J�1m摈��":�ȴ�34���UM��.)Ҡ�^'� `�H$|OP�'�t!�!D
0*w�Ұ8����#��N��u�@X8�?�#�������Qp>��8�(\E�.EBb��0I5��X]vtl���У"�h!1ph�^5!�d �' ���틑|D�c��؂MAazb��I(N~:|Pa�\
K00�C!7E;!�9Fev�hf�U3�~�c���c��O eGzʟ`��R+���`��U�R/
������2�D�D)��������N(%	���5	�&B�i�����{)1O�U���j��}&�\k� �T%� ��7@����C�"D��y��0B��`[���r1h�D"�Is���OD��P  ��Ȉ۵JĥS�x��'�D��F��A-VP��
R� ����II�4.?�	��j1Hdn�0�]�&�Ѹ%H�Л���������%$�M����?����D�3M?���㋁��R%x��̍ccV�2��T
��ɏ��j�� t��g�I&��1�@疧?��e��h�6$qh�Z��^ >��o�^����x�h�hÀ]��M^ X�A2�n�5)�b�D>?�Tß�q�'� �� L̂N�t�R�eZ�3�0
�'�Pt�Bn3m�88"�僈'6�"�&��d\�;A��)�ǟP�'��(1��ǯL�Iɉ
SM���
�3_��nZL�ܜ�Iߟ��'X
ɺw�'��S�-~��u,�Cb�L����V�`[CʁO�>��v��9~�}�FG�m�' ��M�v���`%��*UI�
���H)=<���'dQ�G�I�,�B��LH��E��2�$1X�O8�d<ړ��'����g��8YiU�Μ/n�q	�1��'+�}� GA,�Lm���Iv3�{�睄$��Y�9v�@��Is�X�5�L�*�`���2Lލ��E蟴�'�D�4�'��@�:2-rA�ߊTF�ta�Z�T`X3�'�-1�p�*W%K��Y@Ǔ0�,�Ҋֳo��yC�]�(�p�8�@�<�v�b��κC����w/;O�lښ'}�R�8jn
�H�3oʸG�$���=�	b؞���$��>��dZ�fLB�L���;���HO�S YIH\�FfT6��4���<m"ы�՟��'o�<����+��]j�':�Ӛ�M;Zw���1�%�XMp�狯#�tPA�K�Or�E�-R� '���G�]P@����	�Ev�{�O��t�d�_�}���;��^�	�|�O<A��K'R��m�~��I���iE�j��d��g�\rM���W�''�����?ى�IaӐU[&�R ���������"On��R�D�m��aV��w>f=�Ĥ6ғ��d����'���sJ�u����� %�>h�@��z�H��"�O��䒻\Ѵ�o��?��	���'q"ŪWd*]ƹ�uR& B�}����*�%�F�Q${a>= ��ә~&��#1��){�xhՂ�g����jö%�
���F��aJ�.�3��'Q~=ᆄ�"L�������
�h;��O��Z���i>]EzR�6s�9�b�HK\��M	�y���hp�]�H�S�uZ�\�?)�6O�X���r!�I}2�˷g�	1�A^��|��p�`m�g����I͟P�	hy2���T%B?��q0#IZ�P#~�I�]�6~ )�U4	�z��$[2Q��I;(FtX[�iV�:�����E���3'cJ�"����(���=�edTH�\�3��2�3D��	<�Y��͟�G{b����C~*]��f]�A�H�Zd�W���{�,:��^�hHM#�])�"���J�"M+qO�j e�O(��]�2����Z��o�Lm�
��fo�c�4�$�m��OQp]9�͓3'fF��pf^��q��'�$����]�ea��ET�-T�@ӓ��'��)q�i=
H�1��-E�q��q�'�4���L�`u�W`F�c�ђ���#�S��ݯ!��W�U3�����`��Q�ўs�����'M��'nzi*���C���>+�Fl�y����)���}&���K�x�Rc\Q�V��uJJ��y�Ʌ20��c��ʵ8ٲ�Q䣇�ʘ'ўb>aTJ�7���
P�)�`0D�T�G��<KS�
 Y��%�u�'�哷��' `S���~�:@xqÜ�.Bz�r�'���ɕ!   �   r   Ĵ���	��Z��D	�
?S��8�d�@}"�ײK*<ac�ʄ��I&`�r@xR%`ӎ�mZ�T�Z���EĒL�5�'&K�T��ݴǛ��a���	�d���Kd�N�V&���b� �Ɨ�`�L���	�Iɛ��#`���bc91��;�����NWv@ ��:�	ZV��x׹iz��PZ��I"�P�@�+xhI; ��t#�l`!��kk��	�:v�-B'�	���8�𼪢�Ѣ6߶��6���H҆_�e�֡���J+��F${��q
��_�8���2"g��r�N��xǲ��A [!`�>)�W�2nu:s�@?�ˊS<v)
��_~lʭ���lZ�����9�Z\ e���m��X4n�9Z�Dڅ�OHC��$�Ĝb��4[� r���)D�jMExr�R�'X��' ��w"U!!jF���aЊ].̔0J�p{��I%n�qOJŀ1
N/.D�=��eޗ��3e�i�F=Fx��W�'Z���r�ŌȠ�>t�ɚO���'M�Fx§	C~�b��g¼�2�$ix��W!Ya~Rj�A�'|J1�?�dE1D����n�2c^��( �J�qJ�#<q0�6T8��ϥE�f4���X�Ab���ұ�1OH�����:ˠ�1w��K�LفŎ���Ƶ���#<ɀ�/�IƟ���N���&h�=wT�Ij�ͯ�(�.p��T�'�R���o�[���)��M+Q�v�б�IQ�Ȭ��F̂Sr����Θ��t;*�7(ʓ�~�'���2QY�4d
�[��!I&!]�0�� ��N��O�� �\�+a�-)��,0�@1��"O>���  �xo�ځ�P��y����C��=!��J�	� ���a��y��>@/H�D〟|�hd�����y��� j��R�G��V�!����y2��	��ȁ���t��/8 ��'�P=�@*qq�Q��Al��E��'����ڃ%�(��7	\�Xgx՚
�'Z�Z��,D�����>Tl��c
�'k��J�NƸ�h�2kʝArPe�'�u�d�D1�n�H!�G����'�|ܫeT�#�z�q'!I67w� r�'� ���jR.Hy>\ɦ⚻_� T��'��1��$i�P�!&�T�|�NyH�'/0��'*�v ��C�
�Q��'V� �T�0
�te8��ƛB�� ��'7\� ���2G����؉:��ؙ�'ؘ@"ɬMM���(N��P��'Ibe   >    :IZ@-�nkZ��&C�'ll\�0Oz+��AI��e���X�'iD��  ��م�"}c5@�"O��! /   �	  �  �  Y"  3+   �pA���D���\�'ll\�0BLz+��A	��e�2b������Z���'����3Û�� 8��*� [��i6ȃ�_�հr�'*��F����1-SB�P�Џ�'\x�!���'|���/E�9^��c���2!�r�E�?Q���䓬?�����'w����I#��]`���fHߓ}�'�lq��h7T�	D�W<.��y�{�Ahwr��_�D����03����	�Nd@I�=��'�f�;����'m|�YO~r�E�b8���uCC�0�Ȇ
Ok�<��A�%���F톂?�ؼ�m�]��p�?ɕ��t�����%S>Mm�`x��Fd�<)��Nh�)��<hB�@ �M]`��L����^$6QB�AJ:u���h7�D�y8� ����	2k��<�@��?xeK��0!�a��U	��@E�[^̓7��A��+�3�$D
{�T4����Ju.�#U@�0P!��΁C��EP�j�T`�ER�1O$�=�|�eDCzllV<N-�Lc�.Bq�<Q��U�-�N ȤҝT�q��=�HO�ʧ?�O��:�d�@D��Uh�P���G�'5���;�	�h�v#|rF��3y��I&oPeqX{���b��X0s��K���贀[b�h��WNR��E���)D��3 /�>o�j�	sL�L���)7�#���<i3�-d(�$��N�W!\-�S�TG�<Ic�J�DB���`��<Mv-z7����4�OT�GzBE#�G�/�<�"gk H�i�$J�Up�R�㈋HR�%�	ğ���ퟜȴE_�_�.u�	�|:��i�h�� �h�����[����-����O. ��D�+_�M��RWhRV<���[� �L9�t�F,S���R3��3d��������I��'2��94�����h�
x���"���"r��{�=�$��f�e�W�/�� ���_�F�qOޝ�w�O
�z��T�w���	��0P���ҿ���cWΓ4j�T�O,��ǡܻ^��
�=��!"�ɇ*4퀰����G�>�`�
ayB�K�@�%���D��$DZ����hw(��o?,O�@��'�Y�����{��-���ߦ&����������͟�?��a�Q�MEpIy�G��Y��<	��p� R���\rz�b��c���{ ��z�@����'�?!.O� ��Jpxx�����p~W=K�(�;�@�S|p�Ñj�?8��q�<DrQ��,[�q��O�|��ٶ=�Y��f�/.E*���x@�O��HHi��W�aQ7C��A�5���x�.F��?1����'��'���(ǡ�BMF�قFB�2�Ey��'�v"�`�&R0Rȓ -��~h�2���X�W�X��Yž��C��T `����$5���v��'R�B�'=Ɓ�Y�TB��'5��'q�HߚF�H�Z�%\:�@
�
�Yy�!kF�a<�-��E�47�^��:q� �X͟Vm�O�i �E��!��id�T�su�P���]J=��c,�g2&�ɤ�F��|
u Ŭ)�󎏃�H��P��dá���(��
ٴ�?���n:6���|*���?9���?شb�V���یq�h4z���)�Zp*v�I��8��%��-V����˶4��`!C.�ON��/���M���'|�p�'���2�[�L7����%m��I�2��u�jEY�rt�*.�T�D<>	|X!�` .>��$Q���Y���O����n�	���J�� �/�{���(�!��'-br0:%N�-x [�M�+s�-P`�'���$>' ��C��[�0#��O�{�?��C_�d�&�/{T�`�߶9�qO�utA;���	�q��>OF6M��7X��S@�����R�%�������mkB��	ʟ�#� Z8��s��l�
�ܤ�P�_! �����@�TPf��$^'qg��@v!�:;�nhI��j-[�j��Ў�1uA��p�&��剜y���d�O:Il�⦭Y��-'1�h�3*u@5�ƚ���O6��B≙Z��1�����
��tbӌ�
ajh�D ��T?)YjѴ�h�b	1~:$x�"ԐM��h�IJyRLF�jA4�c�'`�X>ݻ#�Ŧk�ɥtP0����7�*,	�'�*�?I�R�l�a�)"zk,��'���!]�m��!��TT��jQ�՘T�(�%��>4��'���%��?��{Ĭ-kC`y��ꏅW�D�(��۲u�~�&�~!�\��x`M��?I�C(���'��y:ם�Z�&ȸrD��a�T�I*1p�X��^X�D��2r��H`JH�,����/TC�'�i�0	G8�n�V�I�[&�)�� [�r�C�+_8%�2��u�<����?QUn^ln
�����?A��?�6�.� �i�I\%
�1s���<y���c��+r��'�ꩪ���m�܁E{�c�m���X����%+I�|k(}��>y��ێٱ��'oq�Be#%�F����ܰ-s���f�O��$�O�	�r��Oq��I�e�u*�"��1�$�^s	�4�6	M�֐x� _;�:=�e"x���y�i�>�?1#0O��)��I̺!�'��I�)�(�k�득@�P�d	H;Q��R!k40P����?���?��-K�#<�������>]h=p��)�R�(ǉ���J���N���)	�8���;�ȗ* ��X֠Ч?�Ƅi6@P#A�2e���P� �7�S��]3�����{$ϕt�����զ��ٴ�?�+O$�D)���^ʚ�2��:$H���!9.Θ��D�p�R�z���ۀ���j�c���㞘	�dg���'�Y�DX�U2�i�<1��*�
MyTh���(L�Eo�O����M���g��O��ydP���Us�	�h��%�FK�?p���#Ǡ$v���䜒HJ�ȓBʒ��T|��t�m<9�EEBF�ay'�$�?I��?y�4l��BE���-��J�Wf�6M�<A�����O�Tڡ
�*D�`����Ո���0�S�T�O�4�
4�c#Ip� J�W
P6��r��'D剬bܨ�ؓ����8��N���B73՛�Äo�f(��S���E��F�-|~ �d�OYX�"a>�*w��<�S-~d��6(�O�uz񪏇1���ۡnԼٍ���1��'a����B�?Q�����m��<����KJ<5340+��s� �a�hN��M�:��I۟x��4�?�N?��U��&�8���`���`�S�g��"�d�Oj��$�R��Za�"8�Ȥ�P�	�a"=i�OR"�b��n�VO�`�ӂ�_=@M�T��l��	��=���ퟐ�� ={�h�vkڟ0�IL��.z���K߼bO,y���j��q�$׷Y���'�����:T܊]F{��6� �A�Y�e(D(Y���r+��P�>�0�Ľ?ı��'a@��$@��@��0�T"� p��O��D�OD�)�Oq���)����>l�sMζ�����-����x⪜9
t^q9��*2��	�P��?�1O2\6�	���c�'���[mz�R��.#���E��	=����F%�����0扶#�t�R�� ��՛b�i�w�:nÖ(X��I!���x� �ڟuG��d��_<!�$���.��ϛ�s<�@�1��5 B�	���|Z@솿8�R4�PBL�5����D�t�160�R��E��0�t��1i�� Ɉ��ٽQ�u�	"U�V��4�Ov�t��-�� S�'��a���K��'���O~�"%�D�r�"T�t��y����f�<q#��zWj����ʀg��T��(Dd��,�?	�l�t�,��/� *�Ի*�f�<��(&�����	�o.�����c�G����~�� �m�Z1�k (I�i�
8	#�	�C��x�y҈Y8�r�k�z/<�j��y���3N۞ޘ'B�J7��J�g�	+>�h+��ɢI����!
8
�0B�ɈRv���aK��
���O"��c��D{���o���ja�˻<a��{�;�y�*�+U��AL�8	�Ց7/Q�ɑ�x�O���ة�ΤC��YH����t����O| ��cCz�Y�:@E�$$Ћ@U~A�"�1A�	AkǖQM{WŘ4��?A@a�j!�����yP$a�EIv�<��K7Ap�(G4?�9�M�u�'��y҃_<	�h�y�@��nu�d��yb�,I���� ��8��	��?Q�\�ر���s�KNRu���4*�|u2�΀�~���ɘ>@�2D,��>c��Bb@$�D�[W�P�u- a���C/+�!�D�_kz�
D+�H{��i$nԿy�!�D�+\+R�˥+�LX \��hB�	$gG�|[�k��i$Q
:�B��d�t�I9g���r��:�AAgҫ\"~⟈+��*#݀i���=� �����LZ��c���]�l�'�x�A�,����'�>�pM~��D_���@a���_j� �3JL�<�R)��Ukx�J�È9<�8m�XIEaz����G��)���L��E�C녲s^!�۔l8d�҂�*��("DI���O< DzʟR9P��-v
t���jP<���+�\�'nՀ�g)�I�mDz�ɜiP*�aW+&b��dZ�iͨI�Xc����ר-�q�ɧ� �"�b �8���y�f�5V&a�"O�)�&AB�j߆Q �啗�(��� �S�'4g����C4iV>m�jʾO� ��ȓ���ZE-� vf��0���= �S��D�|*���`P<�sЮ۫?&�0��搸'.r�D�xDb�|���"�'q{�a��kD*�-���J\��c#�n&�Ѕ�ɻH�< !j��N4��J7~yBB䉨Pz���!c�X��@�%�("<yϓ5�D����g�"p떈(�x\�ȓL����S��-H<���ck��������{�'��O�Qf�E���E�d��,��9��O�Ez�Ś|(1Onؑf�žQ~�'Y���lDf�`XW ��=�!��'�� 2�d !ĄL�-�>���J��1 *G��IҊֿx��9#� Mh<��a+��������A���
~���l
�J�9��� >������X����I"�N�./V�z���8M+0}���>�A@�q���<y&'�S�S4�h�TA������'��&^�C�ɷ��y`��5�BC`��38P��D3�	x���Q?:J���CCˉ\�|B�I#��p�3	�3����H"-}r������?Us)�Z����ƕ�B_.l 4���HO8Isc$�R�z�8��� [vrxOT.��L�'p��<�6�S9pt��>�O���Ԏ]F)�P��+��Z��(Z�"O�m�f	C�U� Y�g��'�d4�Ş��`"��
 Pk�"�2F �ȓ"7��QT@�(v��M��فf�-[��ķ|����\���Ѥ@.�D��ES�JC�T�W��b�\!��(�'$�lԑ"CM�J�򙉵�5�L���E7)��1��	i-\���N�D�\ђ���4B�I�ff��Ԣ(��i8�Z:� "<!ϓ �6��U+K6/���b8D���5D��r��Q�*�;�Ih`m��(��DSt�'�\�O��� .E��Y�SÓ�qq^�� �Oht`-� ea1O|4��#�%��'�lR���3%����J٬0�lP�'�y³h��~���AdH!�q��'�^��t�Z	�~mt��6%iACO0H����dތBƠ9 <L���'�V�O���a��/�<d�ďE�p�N�Z���B�'�!��"�OXQQ#�OL�����|x<��>���RVv�=�<��d�C��#�L�B�w���P����Pc6B�	�z.}(t�A$ �~Lx��	.$j
��d=�	�e�$�6e̐(�\��Ŭb��C�=���G�A�>�c�_�&����?�1�l�''5J��1��=�|]��ɸ�HO2�ALl�f84�S3j/a׏Ի}�6��3��[vn �<����[f�>�O�i�!P�C��H���_/26N��"O  :gl����	 &l��J���9��D0�S�';��0���	5=����Ut�<�����T4*�@#�T${�:�HO��'{<�O����D��0��J����'�n����>�I�R|j#|��%�B�9���'1���D ����#��R���T��-�((��Y.$bMICN&D�HPFoɣy=�@���2�BM�a�%���<�3�8&��!�q'9n0�aP�J�<�ΉN������DU!�}�ab���<�O�QGz�e%��J
EUR�C'LA�X��i�E¥��$��,8)��d���MkV�7�R�[򔴺f� AI\t�ae�'M�!��O�DI���	�nHމ1�d�$o�!�$��@V���g�L�|+�؅�� +;C�.��!8��I�v��4x2IZ?��@c�I�9�α�D���%,�XH0O�VL㟨D{����Yy��$�!TQ�4�ͷ�B���R�	��l �x33�E�R]r�&?���F�;K+�! �E��� h��5D�� ܴ�2��o��<��k�f)�Q��'��O(L��*Y&���s��X�ܸg"Olp���ק��8�AJI>@ (9bg��E���	ޯK�h$q��t��y%`I9e���Fz��lc�,�����=Y��܌1KP� ��D�!��+#�3�I5ag��;7��|r�V,I�����(AwP��g�#�yR��*;�كNL�aa��c������'ўb>%[C��;jf@�kJ��;�Pj��/D�@�f-��}H��y�P�AׁPd�'�"��'�Ͱ7E��h���dɹ~���k��[l�1O�5I��S&��8���QU�:e��H	/�:��f�������I^��!]�z�)��]�XJ!�҃*e�H@!C/�x����VC�l�牸�h��b���Pb�j��A7&��C䉵�1�JܑsN��I���we��$�s}E?ғh�'�ƨ�Ŧ��.�<��ï}^��'G0y�Ƙ��'�6����� �������s_�%����������
��V�]!NrD�V�:#-����j'f�RE�3e�Qc��3{�DZ�'>��YCnY-	g��c� �U��Xߓq��'dE�_7�L<c�ʵB@��5d>��(�HO�e���Ԣ�İB�b�x��ܹ_!�̫�l(�$c�B���y�@���'T�FaZ� )V��8�F2)\q��8N [�͗�9z����y|�D��|�=����QA	�G3.H�E͒tA
��ȓg�I��I���1�S��zq���?�V�)ja�I!T��1��#[>e0gn��hO�`����j�N��`��y���Å��.aR�`��dK�b4�<�rc�+��>�O�ؤC��8&�H�$8d��P�$"O�y��RA¢jy�Jő@�D2�ŞUE����ET�t���G�H�H���p���K#k'�5!��z��t��D�|��Ē�N�*3��qL���e�C�K�r��L�b���A=�'Q2(�ƪY(S�hp`/ܸ,��H�`F�2n�d���I�-?�	Ha!D�u����%���B��!t
�򔍠7O�7NdN"<�
�/��X�@���@�)$>��ȓFr*LP�O��B?�������$��dXu�'CT�O08��$�Z%�G�A�Ns�4r�O�� �C��O�C�Ms�'������\�+�����H�:��'?LDX��=:�6�k��(�PY��'M�b(�'"GRQ���E�'�*�'O��x6�_#5��X�̖N�j��'>ʓO$X�Q���t�jٺ�O�셡��B�'KxZ��Oԩ!� M	2�ua���]\�1��xҊF�=:.��<��b�{��2�HPχL�hph���'�C�|S00HP�Y�c h��(�>����+��3��`��U�� pQlߤM0�B�I�K-N�I`J��z�
6(�#~�N�$x���?�Qzg�A	��ާ6�4����=�S!�=������$?sx�-�G��4� D�vCׅN�1O E�rKץ����:R���D�
�&��e%ҝ	b��ȓ4�:�Ckم����
���<���	؀G�h��6�B9^�d��Ĉ� �!�^�z�:m���	"����f��"=�)� 9�?�����a��,Q�d!@�͟���cF���'�<�G��L�K�ȊjZ0���)�[m�P�DН��?���B)$@�Y�t"�uBQsBϛ{�<91�JGh�'���|Y���m�'��y�'\(h��kE�Vm��"�y��F&t�0"� ��)!�@�?AW�3��$(扻�n�R���@�����W����_��Y� :�I��u�gU���EzJ��@� &��s%+M�B�h�ȓ?�+���P�@�̚�"O� < �2.D8B��i���x�9��34����� ��sb�&Zʡ��=|O�i$�T�r�V�,��hz�c��a�ҬK�b/�Iz��ug	!�?�&(+pX����S�� i�+��nȚb� h��$����`��'��>~��$��C
�9�!���3MvI��Q)�K���T�az���K�o���!��#Gy�
�`}!򤉏1������h&����0Q�DH���)��R@M��Щ�(�-��]I�퉳�z���yr-��|+=Z0|�ŰZ���F����'����B��s�g�	K��;!nT.Bd�+�탏�hC��%����!
͞9+�<+1�.PDb�<E{��$-�s�z8!	%���b�Y.�y�n�?*���gf
XAv̒�+k��\�Ob�� �EN�x��L��H�<phh��ΉCX��	ӟ��ɿ,�޴�?1��?y�O`xCTB�~�L�A��J�*@!2,7ź1�^��&Ǌ��!(�~&�d
CE�-x�+ѩΨs�BS�V.gV��a!�>���Z u۱��'�p�P0˛�S�m� �TuX�8K�O��$��-�i>aGz���d��	�����t�X��y2�X��9���vsj0	!i��?��2Olh3�����	}�%��(醨�.q�>��FY�ky���
���I̟���{yBe��$!�9�z5�V�ڊ�8����*A���j�هP�v�M�[��[7.7<O֩�%�Q:#��4� ��b%�Ю�e��23�B;tk2���:<O������U��$�e�Z�+�\��v�;/��'WўP�>1*�73jp�Ӧާ\Ȍ$�ׯ�L��|�I>A�Y+6[j��M$sS�Jܓm�!���D=	���O/�v���"��f��r��J�ꑣר���<�"Ջ�?��O�~Tm�9��S'.ɽ<�VX��g�b�	ӑ�Ȇt�z����]8�sgk�=;u��I�-Wxd��#�`ĘQrMK �����ɆZ�x2M��<����DU�k)H}P!J��$,٘���|qOb����9��1��ڬ,�\�ٲ+�GZ�Ov�Gz��0�CS��3(K�%"7`�$qWn��u/�5H��<�%��h�����?Y(�YnZ�+f�ž+����1j�;���2@ÿ"���'��B"2~m�}i4��%�2��O��&@ӟ��C�G|X2` @�Yst4R"�^�IU�4T���9-ʸ�S&EV�O��0W���N��u�`��Dx�%�L<��+�ğ���L�O��6&���1��	Q�Vs�&A��y��
�!��m��ыD��DѢ$G�bۑ��'�� �?!�cQ#GO~�C���7���sI@�`�5p��{�R�'� �kaӼ�)�O���>����-*i5C �� 2mX� �D�	X5�Y��@\�0~t��'�%������3��6k�ڳaH��Ԓ�(��K+�ԂX8wT���1�ڬ�W��x�h� r�H f���;�D]35Ȋ4P���$'?�Vj�ݟ�B�'b�yi�@�/��K��9E {�'����EOw\�]�A�ڄg**��~���
_������4�'3�\�@�P�bȃabH2P���4#ѤR�,EnZȟ�	�d�'0��25�'��i�2&��H AK�
� 1���p�\�Q~x����_K؞`�`�	�0��v�J*<���Q�2Ly �]xzj�� ���LQ��pe�tA��zy)6�
ɟ�Ik�'��OHha��f~�%�� �$Z0kU�'��O��2E��,E�S��*/�$��0��J(R��6�i�]iǬ���&+�	��H8����Na�3�$S���'�N��J~2e ��y�%
GI�&BM��`�I�<�S��l�:M�䇐�2�����C��`�?	Ra�;�|����ԇ�DE
�f�|�<)m�a`@c��?�m��Q��mב��'x��X�*D�/�Z����Ѹ"RP�P��D�R�Y�<AeJa>��d�&jf�xH%������ A̓On�����0�3�� �kU|<�f��!dY��(���s!��2۲�9VgˮFB^�����? 1O^�=�|�'e�n�Abw��#{:ـ�C�`�<�.�N��(Җ�:1������HO��'Z�O
4rsBF5	5B���gQ.jJ�159Od��d�CP 4  �   o   Ĵ���	��Z�D��<&��8�d�@}"�ײK*<ac�ʄ��I&`�r@x2�a��m��>'�t��ȩCL���$�/f~N-X۴lv�6�p�ن�8���1�^�$�b�(Gl�U��_n�'�Dx��Ȧ�"�@�6aZB��
혃f�<�5�@�p])��\~�I�?n�D�o���DJ'N}K�W����FZZɸW�P$-���a�3=�r�͓J�b��ދ���Db>�St����u2g�b�����Tn�i`�� -r��'᪐y�c�0y�d	-O�Tu��,H�5��P�`s��O�$S��4����dB�'��y�b\� ��e0�O�4�a�E�M���L"��C�y�T��ٴu�,�u�{�H����8i�P�bO�$sh���K��V��4�F�3�O<Ƀ��D�����L�Bɱ�mG�'T&QꗀZ�y��OV#<!&6�ɕ*sބ��P�I�䠊�Ctš��4Fo<"<Q�2�T��@
CC�`�>�₣��G�"S�;F"<	w'7?)�-΂?�v"L/���@ eEy�v�'y|��?Q&"� �PԀ"L��K���q���"�#<�V�;xԔ��1��D��@N���L�-Huz��C�O�t�O<���݁�T)d�i�
TX?	�1�`�O�h��&*���U��� ���^�MB"�X>���i`܅p&�-J ��s�-C�"_�����0匏$�&��"M,p &�7?�ZٱSEN�x�Ɇ!ʱB���D&�R^(�A��zۚl��O
8�v�)J54��yFyb�]X�'�t̩��ʍ@0�[&����L9�'5F��@ ��yR���^�F@ʇl? �R@�k�9�yl�6F�
E�U�̸��'�=�y"���b��)pO�l�H�b۴�y�aV.I�����h"�����y��P�v]Z�kA:S�h��wOH��yM��f��8"�E:�RX3�DI��y��&\��	�d"_'Fi<��4@I��y�cK�`��8�S�����5�oΝ�y�mßT�I�g����=Sm��y�m�4F��⠥^1)�c�Bо�y
� 8D�aCA�
vL��u�o��ȧ"O�m��W9��Г' 6��'"O�ę��BN:�z'f�Y�D�(�"O>�� �,~�Hڠd0�"��P"Ol�C���,X4+wɇ	�~B"O\�S��ö
��dPƜ9��"O� ����z)   >    :IZ@-�nkZ��&C�'ll\�0Oz+��AI��e���X�'iD��  ��"OV���Y*q�z �`���   �	  `  t  !  �)   �pA���d���\�'ll\�0BLz+� {�ɔ�e�2b�P�DJ��-���'����cD��y&V�YG�܄+��#�"*D��d�'y�=j�+�R����@�%���j`	�� ��-#��'�֙��Y�&�"��BH,��;2���?�����?1���'r��7CW�z6���O\1f�,�ߓ-��'�4�e���$A���8f�e��{��C1m���$�6;����+}�����G2���ԧ��F�.b��A��d��j8�O���J�(�����U�S2 �ܑ��'V�DJd�A�^L�થ�.y���[ӓ��'Έ}�D��Wm��PU��:��r�'� p���:�7��N�${���+�S��ŉ	V
l�A�U��~�h�ONў�]�)��c� ��w1z�Ha�<|�<Y;�\8sf�-��^<{v�m	��L>�D��+n�i���ͭO�������L�<��(�7�Z�@��� ��J̓�hO1���P�(ğ$�潻��5rwp� "OJ�Z��1R�<�A��9y��c��>�S���\y���Cg�-���`�ёoe"-M�E�b���&�*�'Τ����f�r�Jā�b<�Тè;,�ه�I�O@�����Cw��p_%��C�I�6�s�g�	q�.��傠k˞"<a
�#P\��N�Щ�Ҭ�3w� �ȓd�:a�W�փ w�	���
e���I����X�'`1Oԃ%"Ґj�:|�U��>s������������D������ɐJ��h�Ǆ
ן<�'$�B��smS:t��l��c�x��B�Mg<�a�7=|��e���K��`bB,@�m����=�h�U��~�ֽ
f�;G�Yc�]蟼��ٟ���wyb�'}�O���En�����˼$)NQIf�'���OX�Ö�SODn�	7�N.(�����($�j�$�<��f�c�x8���D,s�OX?Q��<�OS�+M��� �>�����4V�<�O�ÐEκ��'h��XQwխ	Vp��ϖ��-��:aV��7�|�N̕x�\����=CP�1�WFÄ��<�ak��l�	J}2�'P+���r+Y
h���[�D��~��'�b���]*~�8��e�Ǒ?Ϩ�g�Q�,Z�OX8Fz����h��ڢ}�P�A<
��(uȇ�%�$�d�<AHH*��5bS�^I̧E���ݡk������	�h�.�ʅ�J>?���O�;6&�%|~���}2H<A��m��uf���x����}�I�neN#<�~:#��-���(�&@+1-��'$�O�G�'������$��x�H�v��%c���SЎ�(O0���=B�L1�b��K�q*�Ӄ4�#=��O�rP:��,�8 R9�g�z�
��Џ@���s5B�O�d�O��c�,�V J���O"�d�O�}Y�Ԝ9-h�*E_�y&�)�-�,t��Ж�Z5a4<��b�ϕ��ɳ�T�L�������?<�9'�20�%G}~|;��88�rS)N�fS:��%g�$��O4���i�5��C���B�'��&�F3O�V�'W�� '��O#��'"�'���N��&���߁�t����D�; ڢ?�ƠGu��
�|�I���+E5��ۢ$��h�	7�yra��y��P)���F��~ZB��/�}�p^1 }��Y&g��U��\�C`��O���<�8�u�i��@��y'�;ZP}��)V~<��r�<qd� 07�D��$O�/������q��6��O��J�-#�V��6���L���E�zP0�Q�\�r��2�l� ��	��qX��Hd��\:��!bc�j�V��=IF�5��,,�@Vm��<��4%��lc�E�'0�FI[%�5O�yPR�'Lr˔�q�2e���'���ȿ�X����yR�iO�0z��R���8�!�?l�<ܫ�{�vM�R#�;L�^��ā�O����+��D�	h�:��'*T0����?1f�iś�͝�b h@�e6�
��ӵS����?Y��O��'LʑAd�E�`!��߼_�`����=�S�#��8i�$�Z��%`� ��(�!����L�z�6Dn��0���4��M����y�څ v�2N����	�]���'F\�Z����T���O���xX�-A��'}
�	cW�m6��ёv�#H<�q�׺��"g�pt��ꀼX�'>�#3Ć�6��$�iL�z�Ľ�V�(�d��	���'h�6��O��OD�ͭ�b�B��k_�^�򘫑f x��D�=��Ӱ<�V�4p���P�G]*E����J�)�hO�i�2�T�o�~�	�G�HIP@��0�r��S"[�?���JtX��	̟|j���7��O����O�S�? ��#g��]q㕁7�`��#A�J�'<�тe˙}��E{�/�/�1J�!
�:���1���6��aQ�>Qw��#yM���'}ƍ���/�v��p.ݲ8׈�h�g�O��$�O�)�Ӎ�Oq��I������'�V�㮃�aN
M�M�(��xr�4G���2�0ї/�+8��iR�'�&}��$�;zxY��ёIϳ ����t�ib�S C�!���+0�i�B�':25OD��� �l��5��!Hb�;~�9�ϺR�����X����� M �a|Ri�}|&5���I����E�6a<`p�!��S���(���P��4A��"��BA��`��8�4tś��'��	�� �>���ǡ'_�@�2��-Mp�!�A�D{�4&��@ə
�1h@Թh4��ĭ;e���	eyҨ�a(����'(�f�.
`A��X��LP��
�5nH�Y���D-xˢ�$h>)y�+�:Z�$[��h5�"QgV��	m�Q�b�8,OhK��B�;�v�/O8�y����~�>XЗA�z� @���'�&���?A���M�GG[�2�$g����B�H8{r�	ߟ��?���^:�`����[Pig��t�'�ў�� @�H+u�ܘK|��p���=,�x-I!����D�';J A�eӰ�d�O�ʧ,�E��4e�F��t�i���3b�&a�R���'b�QZ��UL���r>eӄ.� =���_�z�YǎD��uD���ē?\�$	ujs������Lt�!~�T�9��L�$P���R.2�'&R<{��?��iE��~�Gh}�}nT�H��r�X�d�a�	2���Ԅ剩27z����r��t|�($F{�O+�\�C�c� Ozu�TF�gBPmS��� W�H��$�����O���X��u�i#B�'bB]��!�$;Њh�Cdã:��]�)f�O������!%����ϣN��т�i�S-�jצ^)G�^��g�3}⫀�k��c?O��S�Hߎ~b�Y����"�@a����Iܟ`"ҎƟ�>��M�����~�
t�deʈ3�"8s&h�h!�˓@	��cǧ\:>
E���2E�$y�X� 6�u��Ot�G�LX�ȏ)f#��{���6ӎ��'GL5��� D�'4�$����@���*���G��D]�F$<D������xł���	J$C�,1�
5D����\�*��A��↕18a��
TPh<�Da^0z�<��tl��XG�4�&��g�,&�
�,ȏvW�XhFc >|��ܣ!+0�O�5���'��RC�Q�܊��`��$���*�}�	k�n����mY�g׆h͞�c� ±M.x�RC"O�r��>!����y  �A�'��OmH�)R<Qv�!��/��_p�`�"O����aD�R���@e���J�ͫS��o����ђw~�K��=��s�C̾�Q�Ђ�>�	D2R��"�40�!��O�D8#����'2"`1�3�B�<Y``�y�d	��Iv!�d��P$  ��)��DNnt�OQ{1O�=�|�tI�j�4�a����J|�6I�@�<��j�7L3�i�E�=���ծ�;�hO���`a��C�cC2���UK�,�FT���iڌ{R��(�V��6l�EA�'V�fn���w��I�d�9��v�pL���%$��90��:(�p���2ū��")-���elA�I~��Dx��'���)�KQ(���cSꖽfN�
�'t(R�,�tJS�W<+h�4��'F�	w��0q4�S�S��a���$#�L��A�>	�4r�b�Ey�/�I�hw���,�V,QW'ڦ �dC䉲{^��w��/&:D1 �/?�XC�ɜ�}�0�׷HP���f�:�Ɠi�zy�D/�5h��E
�̔!xG�H��	Z�	!ƀ��C
�2!����e阘n����D�H{2�ڰ�����*S�28�0FM����'E�u�=!W&.�i�d<,� ����B����	`R!��P���&t�hqR!
��N6az���n�h-y7&�b�h2i�6.!�Q�&�� M(_�jH���]�Jo��F{*�̠!�c]�6Z���\�rبp��%�W�'�8m8FA,�S�?�b� 8�r!��/��R�K)D�� ���'������,@<L`r"O�41�c�
�fx1�劍T�Iir"Oj��4ppЈZ'��$-��"�"O�-�H��`���G#L��2�if"O�,!G�,bҬ���aU L�ڌЇ�O��h��)ڧ$�^<� ��=c�"�T�pC:e��+��e0q�A��Hy���8@o&���<�ډI�a���T�ȥ�2���ȓ,HHd��õSl!(�g]�^B$��:"��qE�B�����Q+���ȓ��46C�#ðÑIxԤO���q�'��}��
��dl$�)�U��	�'���Q ¥����'O�4o�9��':��6M�4Jpq�ǉ�Uw���
�'�${V�p��h���HN�$C
�'h�
���.[&}���!>�����[��\�	NF8ì�00*���#"Z))o�B䉿e�Q����n����`	�B�ɕ%T�"ե7&�>Mr��"J�B�I%� 
D�P?q�C�)0_�tB��	ҠԭC�؃W�*g�B䉡>
|@	P�&Cz�Q`k�m*�>T/�k�O�L!p��H�J�t0�χ*{�>���'y>�b'��w&, �&��ٰ"O���kZ�rZ:�[�@^�jk��5"Or��.E.s<,���͛g���BS"O�b(�������K�M��"O���'H@��,�Ʌ&7�r���OL{��)ڧ|�D8T�D��U�U�w�>A��gM\}���ýM��p������ȓd�<TZ��E6�iAp� $�F�Gx��'bE��R�+"|X��B$93��J�'A�a �I�p@��0��
2�!Z��NO�	 �HOLb�����A�n�����/ q��tH�䡟�+ش"��GyrBI~�	���H֘T����LR�l��C䉡{b�]Y�	�/k�ȚD�J�O��C�ɪ4b�8����q��\#1T6f����)(��3Q�̝@�
u*�!(X ���'��]����cۮ b�e��cX�x����?����(0PF�'���c$K],x��D�Īf8�҉}��_p��RL$?� �N�:��`9�^Q"#�?D��j$Ϛ
JOh��/�Z���Z�d8LO��ds��;#ƌ�w��;�b)�g�:D��y�/�ok�M9��K�>s���"L5�	��HO�.�eq�@�:���1��W.nF�D{��<�bc��ڥ7�^}r���qb9:�D�]��M��J=��<i��L*v��|2e�8F�ZLX#��(�T٨G�/�y�hR@����d�&��Y�2/]�Ҙ'�ўb>��`-70�!��^?l�Hd�h>D�����ܒ]���aFM�"$���aP��E�'��S��'U��`&&How����Ɗ_�\���Cb|���L��(����:��g	�%����`ϢKڨ�bQ�'��A�ə ���r�Z��5k�'�@`c��ߘ�
��f\	�@Q��-<O0�(�%��a��X��ڙ�m�"O��H��=���J��I�\��CS�'�����,�<!e&5���Q�קKhL���b?!��i
��A��d)���4!Mܞr`8��O1~�6���>2�	&w\�b�L3?�X�ȓL5�y�G�	S6<ܨ�!Q�r��Y��'f-�GD�:olB������a&�I�(��'���0��(?t5߼{�Y2��)�ӺK��	ڟ�g�֣�\�;���>�L�75�I-H}1OD Ɣ�$+^$���	��E�%ԍ�X�����S�? z�*��� tN!@�=|��'G�OܪҬ�^��Ơ��@�ܕ@ "ORM+@E�{���/J�M��U����]H���IҖ~6x��
Q�lǼ�������=y�E@�a�1O�`y�OH����,m��YJ�K�"��q���"R��MA��L>9�
!u�a�`MWOc�gn�<i����vbn��!ZuF,<��j��hO1��S䃗%b��%�b uw�0�6"O���s�X&:��#B���PA*C�0���^z���U�7bV۶N�0��@�y����IܘHڋy�bTM��?i��mɮ�Y�M@�	�&}0S�K�c�J��
�6}J:7,%�egۉ*�M�7��u�<��S���+E��E�m��k p�'�y�n�@�HA�U�6l@ʱǑ�y�mҀy�~Ҵ�����
w���I2��āb�'F1O��EJ"7�H\�T�?V5$���O��m
0:Ң<�A2��Ȱ98v�aGT	}�ް�RD��4�!�$�M��mh��7 ���Q�	P!�DO�_�e�fI�#D�]ct%�PIvC�	�1��Ι9�R`�'L�Ffv���f�	S �ղ�%�!Y��r�R	P; �$E{Zw_���jN0%p�R�u3n��c��<d���>1�� �� /a ����0u�օ:�z���7&6<� �"OX�i�ilEe��{,��'��O�Z5)
 g�HZ�/P)Ng��K�"O,�*�ϧ9Ĵ� 6L
�|Z��D^b���	ޅSF�P����^��4@�k��[wN�=awK�Qk1O�<a�OI����&	#� ��'\?ِ2v�d�&SR�\���L>���ܦܠY�'ҟ6Ϙ��i�<!&'�N�`���ߥ�N!(G\h��hO1�`�0s`�F�݃Bi���t�q"O�`��#\A��)J�	�* (��8����b���Q)j!p���2�o���	�"^x���y�e��?I�k�"yB�@Ɇ��|Њ��Ǐ�Y�����^�h�m��YY!c�0��ȓ<�@q����	C-�Q1CH^�s\&eEx�'���0���)A2�R�!}��eO�Y�<y�n�:+��Q�j��.�Dd��)[�<��O\�Ez2�dñ�]Y$O��#��@Ӡ�,)�d��:�����f��'0�m�'KZ;W_h���C�SIr���'�2����C;$(�����L�h�k�'7.�ᣖ><�H���;pf���O�xC,I�&�(�Ӳ��s���R�'B�O�y�B�U�,��b� q!���D�i�'�D�+!�O���H�z99Ǩ� �UP�>�A��R�8��<�p��G�S�)�p�P��5đ�L���C��&�.-�QJ[�%SXy�/b����� �	�SL:�:���<8Ij �U�Ji�C�ɉ%�����̖!q�ʔ�va�
G��⟤����?-Y�iY W� =�2BX�(�fyK!�P�'օ��'*�ID�Iޏ6o&as�מ<H2���4�.b���0���q��'�������B%Ҙ��-_nn&̪�'c��hE��`8�a��ɇ�1u
캉y�)�S^�jfI�3V�ɳȉ�~'nB�ɰz�li�*�`����' ��f�R�Fz�[>u��*g���P#�S/HFm�%�Y��?�°J�1O�����'"��x2([%>�r+�NϚU��Pv�J����O5���"��������y�"��lv���ŋ_,<M q���O��$]�!xG?hٰ�i��̗k�!��]#O�tA0	�.��ջ&[��"��>ɑ�	<���ډu�"C2ܺR C�d@��z8����(O~ RM>��Y܆���,$�-! �^�<��s{Ĵ0G�C���t�.��<� ���@Ɉx�	��	����P�,4�@�6���j*����S����$|O�%��")	O�hm�c#٧C��
4�&�I��HO���dJҦO�H���Hċ*R����V���'�xl�<!�b�Sn��e�܇z���a���9hC�/r;q���Nr҆@��NP�kN��$ �	�Bδ��'���w9Z��r��[U
C�I"�
�(�Y(LD ԉ)F�`Z���?�(�@�$��Trw�Z7Tݡa�Р�HO���Wb�m�n��'O�U���?{�L8�@��j��)�<�f��j,�>�ONe�8jT�Z�	�)zT�Mr�<)f%إU @*VoZ�&�P�@#�Zp̓�hO1�xx:�ɍ	|`��:.C8{N���*Ol]�gBO� ��A��8z9�T�Ik��*�	�fMИ3F 0��Z�J-)�z�D����	�f	��M���?Y����d/u�x\z�m^�>����1��h�H���p���.�2�bçשH��g�I	w�4 �c�(��lX��*�)A4� '[�Ɏ*l��X��L<�@��>  �ikv.ڨ|��7���"����q��O�� ғr�LK�/�/c�`��Pj��&X����$�X)�.�8"v��R��
T9����y���O�4��O��U��Ku�	;!�D�3/ÊJ�0�Pc[�K�l7-�O��D�O@�t.Ek����Hǹi� ���d��E�t� L�e	�M= ,h�ǗG�yb�A���8D
�+�^AW��F4�u�C�t�0���m�C��y2����i��A msT��,P5�U����?Y��=�I>*ph���z�6� ��3_�.��dGu�ɘ	+\�)�a���ܔ#��2*�pj�h���,�'�V$Љ�~ڴ\l��"���x��c�C8�*�E�'��
O;�I�	�|:�Єt��L˹<�2ep���Q��-�3IN�;a 8&��+xiN��D?�0< �&�� �88 a��Kz��c[�r�^��D����}�
�n���П��'&<xg�ŭU�� ����5G�4;�{��'�̻��C��x���ѥ(�X����<�S�ċ�?�5 �OP:Gj8�ׁ �6�NE(��'��	�:��H:5���v��	Q��k�^�]2X�F�9��F
y�/�,�4�Ӫn��hCe�~���@2�?���s>d�#���5����$䀫���&,"l4�C�xRl�y7�XA��%T�.�����{�x4S�	P�C�����AL�O�|9T�'�R���	�������t�T�c?(L���(D�d��o88�*]�FU�R���Z�'��	��.��O�}�2���~�Un/D{x`��O\�+�x�2����	�E^�%�ݴ�Z��?�O�Q�1'g���L#��`:0,�.��{�K]�?�pG<4�U�4�L<�AGN�n��T��w"��Aڱ(T�d�xK��$�5kwz��~&���C��q��j�bĩw��	x�b�8�?��O2������	0bX%��@�
$dSD�/M��B�ɂga>��S��e��] !�
θ�DA�<���N���0�'�ɻ);���끠D��ZD��8H���' 
X����?���?���6D���������P��L���v�=J�̚ g�t�Ƽ;�$a�<lO�}a�ĉ<R�<�;����%��R���l'Bp"��1U�d�퉉O�rI��K�/Gc����n�*M���7��O �+���'`�\��ޖ�.��$���BC�,hߓA~�'�P���-�<�ZՓ�!�1c����{bo|������S?=l�#+�t&�S���"���'4:Q�$�''�*O~R5
ʐ=B<Y�e"L�<��b�ȓ^�<��ϊ�}��a�Ê�] ĺ�i�Z��@�?�� f���QCK�BԒ��aJ\�<���4r|�{0���Fi���U�G8���'%��YP'+
�@�"�#���I��q�Ɉa�Uh�y�&����!�'X��Чg.�e"����'8X)J��H�g��ؒ�)�2_X��PdS�0�FB�ɇS2�E*$��&���E�з+��c��F{��4@� I�]+�E�.K0Ȱ�B���y�'݁xz��0��C�;lp�A�Ϟ)o(�O�����#�CLܼ⡦��@�r�٦Ku�p���{��h   �   t   Ĵ���	��Z�D)E�?,��8�d�@}"�ײK*<ac�ʄ��I&`�r@x�Gn�x�m��c�$��	ڈ|��E���P�tpش�vN�*I��I!����ˈP�$�Ƣ�)B�R:�,/�=�l"<��c�b��a�/<�"!p�M:8�Y�P�h�T,��4��PG 7?�5�.w��7��C}��	
�:E#�%�a1V� ��-yF�����4]����@��<�D#�!��A��e�O*擞G���`*�'SJ h7	�wf�1f�I�M4H��T�8x&F�!%���8@˥<��'G�r�I�#'���W��%�^ّi˚z;xd��'������[Μ�O�l	�g���MK���G�T�uź���'Ɨy�(�bUI~��Y���5�lٲ!����4�Y#�<�U�D��O����������r�.Pq�Z�}2�,s��Q��5��#<y�� �I�r|�
C��z4n�5K�x7�Q�O�5���D79�q�ѧҤp������}A�c���@��O���O����"]`(�W%>D���S���Q�.Q��O*M���;_*�|�dAO�$|H�Bʹ�O��a���Z��?�����<���ݍACV�ɶ��H�>C�#<AƇ7�� A��`a�H�p6@u�r�7����Ov��K<!!�'yN-ɠ�	vAFC��Z�����T)�p�l)zߴv����ַ%�$� P�-��q�p�\�*t�B$K�3o��V�K&m�p+�����e�����V���ɫ2V� �&�8�V�Qte��h<�R$�8o�N�<	�	+�JӶ�*���R�(ԘčնD|�e��_�  @�?�-�|�*�<29�d\0!���`��[r_�x�B�N�(�Å�)┨����0���!@(����?1���?)������L��.�OB�Z$J������En�`�t�0lZ��p�5.?�RP�p��������+D3�	�~�>�����H�x=is!��z �T`b�`����,��*���,��$�=� >�0%�&GG>X V��2��y�W���z���xC�O���Op����{p���S�$(�+��a�=���۰2�6�d�O$���E�����=�"���ڦ��!p���+l.����1l��T�.M��F��V
���$�܂�4�}y�iq��r���<ye�%	~!s�̔$!���vV���P�w��@
�lyr��Od   >    :IZ@-�nkZ��&C�'ll\�0Oz+��AI��e���X�'iD��  ���� ���X<�t)�%Z�O�   �	  ]  \  !  �)   �pA���d���\�'ll\�0BLz+��AI��e�2�=yH�����25"^��j�A ��أ?�d�R�IUx��1�J�KM�Pq�́�8�\m���?�td��@Ix�t��̇��`S�A�A�D�K�,Ѯ���$�OF�O��d�Onb�؋w����j�0�N��_i2�!�(#D�t#��-����+5Z�A�'�3��q����T�	���'+��m�� ����Z�(��H����O�5 �KъJ��O���<@ GҙW��o!$��d"Ob�k�LH����b�ȝ=C�~u��'s�O����>�j�)���:��$x�"OԉJ�b��4ӁY9��a��D�d���i�pi�9)C�N&�
��2�R-}J�=aA˃��1O��a�O�I�NB/?z}� V�ud�@X��$
qm�d��L>q�[�+t&���Y�_T�(u�\�<�"�*�� Zb����n̓�hO1�@mJ�&�`'�	�n��mw�@��"O.!�c�2��=��g�>_�h�O3ғ��	s���-�R���E\��JP�~|I�	/j4a�yb,A��?�g�.A]J���H�}�9	W@�?=q��j��	��,��NԔMH2�O����@
�e�eG܆0�`�ȣ`E� Dxb�'�v��B�*2�B �O|0�5�'�޼K�ȍ�x��(��o�`���,��I=�HO�c���BB2������m�tP�AF_<n����"H-�?���?a�'����?��O�&�k"*H�z�:�k1N�;	p���#�x�D2WtXˢ �H���$�K�o���J�'Vvh��Oܢ&�����V�?jV���O��?)���?������ONc�t
RJԄ/�F)ɶ��-L���g5|O^&��1���<�����$��1����`�7�	�9Ƥa��hy�#X�y��3�Q?r6DV#WPMk��ϤrJy�u�4񤛟C�t��I�T��Pk�O�06 Q�[!F0�$�^T�	H˓ !a&�d�$��5�!��6�{dk��ay2���?����D�N�,� ��i�%Ҥ��e����OT�d0�)��3m��La�j��P���O�� �����T?�x�%�D�^�Ѓ�7SX�aܷ��	My��ܽf�6hȆ���Oż\�;t>�Rc��z0�ä�|h��L��!��1}x�(����x���a؞�wlεM�z�F����ēB�[Dx��$�H���ZT�C/z��}�V����_�D����0$?�'>�@F���\�%��T��	zf.ʓ�<9�Hvs��㧛�h`�5,�HO�#N����bcѰvJ�`�31vTd!V��77�X3���?q��J9��
r�԰�?��?)��-�`=����~�x�ED٨v��03�dN(z�.#�@�>id1ԫA+@+�8��Jj��.9}���`]]@�]*P+�&8>�	��ݍfn]�v�L=I���@7擤{���j�w�5��S�)�@�(����R�Ӧy��ȟ�P� ���������������Vk�|��Yp�N�-���S2Ʉ<��Or�!���KR���(� ��,�U���G�c#ң~��1%|����M4?�D���OJ����MKe�V��p�ܧ��áĝ��~���4�I-6曶*�U����F ڐ��{n�Kf/J6\�("Oȼ� ��3�֤-@5g���A�=�!�D$0令S�![�%bH�RE������˳�'�����։-b	�q�ҝk�t���ޢz�{�,��=�PIR��̑l���f�I$WqO��ld�I	�z�q�O"6�7Uv�)��Q;rY8�C�*�0	��	\y.A*|{"�'a)X�Њ���'���LɛK0��A�D��,>�Y������<�Y4J�Y�A�X,�U!��'@�*�G�I|�@��%P'A���	˓����I��8޴�M���PB͆�
�CG��k����^���	Y��|�K<A)	�lLԠ�畯I�&2J�'Fў��.Ȍ�SwHܳ`dؘ�W�q�DP���ȟ�'�>��bއ")R�'������l�
F�@�aB�G:e�L�2ɗ�G�N���?�aC/�<��G.S~�3�(����	�?�Go֔.�(�y�m �px�b�j�	4P�x����&l�*]�1�չ`��#�-�_!�T(��+Ơ�bn]�;��'	T�)���?I��i�~��Oj�� A���^��eᒇ �d:���`�2���,��ɛFxt��ſ\g�h�U�h� �E{�OF��l�Or���5(��,��T�v� U�A|�ٟ|�I�T��p�X���O��${��=� ��)3M��} ���+U/P�((�k���'�4��w �9d��E{RQ�M���Y�Rm�G�֝�z��>Api�����'X����R	id��R% L"N���P��O��D�O� ���Oq��Ȧ�A1o '5L�P8�41������x��!S��@�KO�zi3$bN��y5ONy�$�Һ��'��3B8�z6�>��j�й&�<9��`�e1�&�'���'��K��I�|"�&��
r!��K�rrl
�lp�E�u�ؑ 0di�f7�O�9 � (q�Н�焊��2� h��4��H+�YO9a|"fZ�0������ e�l|��R0Q��8��5��Fiu����<)���'�l�C��^�'���ϘH�(0���sLEz ��
x����\��MB�{2&�V?�,O��P-ƺ���M �Y���8�!��60�!�GM��:On�a�C�gv�1�2��&�:L�e -O����A�*��\ssf޸(F�H��'P�(��(J>h@�'p	q)�D��d�R$<���9�/�]�Iԟ�����9Ζ��`��� H�>�Nܓ�����D�O���?��w����ĔlAf8;E�*��hO�)�X9���W�Ѵ4�L	E�#C*H��O����)0�i�r�'��Ӂ`>v o�<6:X|���=��Y�Y1Vy����?m��+�m���Dm>�bf���bO�32����)�	"z�
1M����:d�lA�/_&Q� \.E16�IR'�S�Sd�4��/_�0�&���{V�O�Ih�'�B�b�l��,�4�����G� cX�
���K�8@���Qܓ�?�
�3�V��Tn�8�{�ƻ6L�=ڋ�ԟ4D�C ���&�8����f���4M�3HցZW���L.�IΟ���D�뮁#?�2�'�1O8�Gʁ�fHM!Ea�k�9 �8@҈ �K�T2�F� a�J��E�	/(ࠡ�S#���p6��lu��;�Hc��4�|�~&�t�c"��8p�Bm�%"%^(��_��?���?B���?�}�'q��I�Z��Ҭ7x�HL�%L�a�C�	�"0�9WK߈[���[�b��2\
�I�<A�v�'����\�'L2��FC@��ҨbAЇRs��B�O:7�R�i{Q��v�|b(�)D��eHa�̅]�DE����!�y�Ľ/P6x�s��jr����-G��y�	����lإ+��[U�(cc�ǩC���Z�i��da0���n���:�B���a|��|�	)�p�Jp��;Th="�F&�0?��̌�?���Q,y>R��S�M�a]�0 ��Wz≛��a`��K
��'O�R}۱؊b��U@b��`'ՄȓU�"L�� >=	d�@��F+rЄ�IR�#S�=� eľP LP�D\+p��x��X�V�Kw��~0�p�ǝ)XMTDx��)j'����}�Qi��4hZ����[r�'D|��{rޟP%k#'O#�,���V.)�̤�2G^R���L<�C �L@��\�D.P�,l�<Y$�ό�^��#E3_g�0�cE�R̓�hO1�h�� �����+eKX�jp8c"O��Y3#̖�5�$�<MY� a�:�S�D�[��.�hBAR&��vF��^E�$7Y���l:��}1��3'Լa�
G�Ю)��CF�����<#<:QRm-RP �-G�+�C�	�Svb�qk�M��Q�ŜJIT#<y
ϓg��I	�FJ�S�� �����LR���Rj�u�,�xtRVI[ń�ϓ��>|O~!�Do�`����F��o��Dq�]� b���J]qO
��U�����P����#}�4p�����gr@A��Gz�����R0���N���~o�p�jͭc�%Y�\&Ӝ���'�����0�*�k���T�\��	���(�^��v`�/G���X��;r'$�Op!���'D.��3&�/X�p�e��7��@�}2��wܓ?N.��TPȗ+��R[L���ԺP]\l6D�<z���7|��P�Љ׮/|<s��7LO��p�K�:P�h���+V.eK'�4D��8�%�*����֤ԾJ�>,H�b4��hO���Fe�"a��,9�Fֻy�>�ր�Y���	J�#x>�@�Ͼy������5�qO��)��Z�g�)� �Ab`͏j\ҁ��MF%f`=�"O
�@��R{��􋇗K�h4�a�.�Ş �%�p�K�3B4\Iu�?T�q�ȓN��}`6�U�@�����UKr�����?!�?��G�UQ��UXdgIYc@ }?q�Wܓ�h��6$IcXơ��gI��z����
�`1�'4��J�bߘM���Kp�T�|ZD�	�'�^�#�X��|z�π?h$ш��.<O���\` 8v��n�C�"O�$K�.�.'�n+�Gþ/YJ ��"O��Ԇ��j�D�Q�H��m��5�c�>�T'N]�����>�Dy���4� �3��;D���� Vi�D	�-C7uFP��9D��7(I� ��m#�f�?Q��Ɂ�9D�t����4+	0��Պ=&�JƮ5D�t��I�
<���C@7t�hxA%G1�O�4�#�'_� �bj1K�|@1ʞ�z�@q�'e�	"#�:|�ȁC���Hm�
�'��3򍎍L��	t�ʞH],��	�'�40*V���zxYA�$Ȗ>�H��'�څ�� Q8vT���&iҨ$��9��'g���&ܿSXМ�&�
q�ذ����#n��>�Ł!S��=ч��/M$v�� D�H��C�bZ�E���Fd]�"�*D����iT�7�x�q'ŸD2���(D� �)�Kv��づ�e�L���&D�4�����&����`y�A#T�d ��5��CS@� R��Q���OP\s�)�'F���aG�Y��dȻFiT�Xk�p�ȓ 
-A�ӥ�i+�o�,������mz5j�<M[���T���j?d��Z�h7�H�ip��|��RԲ0�D�7ef�zG�_IٺM�ȓL�A��J_ z�	w��UT��O�	a��'{�,��I4%�*D@�a�/��A�'�-��%YT
�CS}�����'��tq#��?��=���ӍX��'�h�2�VJ�t�Y �ԡx� d 	�' D�Aģ:]���D�d��L�Ml�}�I�H��Y��!ɭw��eǘ�/��C�	Y�v�He��v���ቚ4�C�ɿp����Ƈ5l��rU
�'F����9�IC����OV8Q�^�3��J)�B䉝�B��$�AP�f���B~:�⟈i���?����Fh�Z�(Ջڜ�S�XS�'�j]��>扡����E�DpzQN-M=[�G�d:.b�����$�q��'-H٪t
Ϫ~�9	���i��q��'�p��I�$5֔(z�� y�u3�y"�)��%l�Q�-�
H��mq0�(K�\B�-[,�������6�dȩ���B�<Ez"S>�@�2��T����*P�h\v(��?aA@4ET1O6����'��):Q`0Kq�p �)"	��$�@�Z���r�بyj�x��J	p.|4����yR�1iqs�=c��!EA�O����|FY�ET��@n�?!�$�<�jeYF*��*�2�b�]]D�>�5��q�8�Q�'C6��� ��674��O����E��(O<H�K>9��7G�2�oK�^����DD�d�<g��C�|!������msql]�<�vH\�DF����͊s̈;c ���x�ңnS���W��- 4�������=���|�n� R�!SF!����3EM���'�ў�]%1X(���G���fc�y�������OPТ�y��ߞ���v���JؼP�)i���:pň���S�? �sէ�:��M)�,P�9������'n�O��R��pBj����R�H͆��W"OB�4Γ�R�2��"St�� �v��HW����ηJ�(1x��ԈP��%��(X�:�ܢ=��M�5�1O�(O�,�k�A�-R�f��$ж0%�����D��]���b��L>)Ӈ�{���!⮊�:�f!ʑ�HE�<Q�F9@�a����
5�t��L�H̓�hO1��U)#-&!����þ6°��c"O`�٤+P�iq�0��� �P���(ғ��)V|��OG�I:��'!����aOO")�N��	�sGr��y��x�O������m��M�7�L��h�x�v��I���'�\�󄀦�=8�m�<����'�����L��)�/ҭ�\���d,<O㐌р}뺅�cG*N+PP�"O~�P'��qr@aQsݼ9<r��b�'e$�XT���<YnW�8�Qs�.*�8"��S?y�i�r,[�y9OfM#I>�Є��[���3&���+;v���E�<A�/Ŀb5~A��+��z�Xh�`DE�<�G�0:z�I�H
�d��X%�H'��x���5q�E��\����� ���=s�|��!�AB'�'v,���Ƌ7��'�ў�]�{���"F������=�bM��Al��y)Z@̓:
4'?	�  A� �d���"_��\�Ѣ"/D�x��]g����t�G�J��hc�-LO㟬�B��$�H����J��af�&D�+��Y�#Ā�HQ@�*8�t�a#�ɏ�HO�>g��t���_�t��A	U">'�%D{��قX� b��h�>�2d���EYۚ�b�c�/WJY&)*�		:zFX���|҃��2�13r�G��vi�����y2
��Mi\�[�GӅ;��L(��G��'�ўb>9�5����b�۷��3?๢��&D����(�4{��b��:u߾����W[�'x��/��'ޔ�� �	gi���4��o(����A	�d�a�d�(��7�S�v�Νڇ���8�{w�%Gq���R6�O�i��G�0C����P�8¼uC"O��+�)o�����E���4�hx��8Ef�BMpH��Mhd�rF&D��@� �b�(M��M�<��`�wa�O��'�v#=a�yb(�V|���T�$��S����~bӴh�u��a�kӟ|�.�$�������P���2B	��y��_cJ���9H��<`QKݰ�y��"�@(��T&s��YyP����DC�r.�d7�X���O
;��{R�7�$G3[[���)�;0�-�EA�G��OĢ=��/p���-'~�g ���%���$W��w����'<��#L~�h�f����Q
ͪ0��GE�<�E�P+(�	[F�~�<dk!H�v����?93c�VE���暴P�R,��W�<�� h���B늇v�P50�/�T��0P���1+�Ikb�L&T���#؅8�	�i
Z�J�y%K/��&+¶B����쓠	��8!PM���'5HĻPM�@�g�I3ET�x� �7/��9���x�C�I�\����!g�>
s�I�b��b�$F{��4��1?�b�W��r���
��^9�y@
��h
p��?n�2q8��_����O�����ڝI��E�D#Y2W�=�d��O�acƅ{̓[��eE��D30Z�v�`��T�fN�*%�ڝ� ����?ad���O�"�A���F��qNYX�<����DL�����
u�x]q3�]�'�yRe� XÈ	�t�/s��!Ӑ�y"��Ny� 0�P�N�ʱ@э�?�V�����?�ɛ1�K�1=����E�3����M+�@R�*4�(t B�I4�}��î�uh�ć�3K�B�:f��Q `&��u���7��w��B�)�   �ӫQ�p;T�R�scL)4� 6�щ�v�3լԒ56�!K�	5|O�}'�P�$�E�(v2����.����s�I��HOD�{��ʟ�A�SZ�4���>]`����3�I�+�1O�L8$��īŒ)o�!��(W><�����A��y2�3=��e�7,W��>�:T�մ�0=!�b�� �L���B<tA3����y�G�+4A�rꃰo��be�3��'^x#=�O�D�iQ���Ai��>U�RB�)ғ?"ISr��J��y'dU+hm��`�Aգ&�\k��	�r:1O8��R�������F��^�\�nT�@�4/0�ȓ%��HX�R�ds���H�H�<9�����-iX ��E�*G߈�j/�;�!�L��� ����\��ȡu�'n��#=�.����?)�EE:������)*li�3㏣4^V�'C��'��+�lc�*�$�O����Or7�ճ9�h� ��P@�5��Ȼ:���L�9#���3i�&��p��g�+���A�l��G�r����/�P9��o�����@j�uyf��x�I�Nd��F�Da�����a�P�0?� �����m�'z�	�hւ,P�#P)<�I�'OP�;S�A52����0�Z�
k4�X�j��7���	��T�'&LB��W7kڈ]@�ˁ���;T��0��hl����IןP�	ǟK��̟��'l���9\h����$���G�(�,���Z�Ex	ϓ zn�����IZ�U!��-����a>��u�����
��	ϓ=��ٸ�/�^��-ۗ	�Y��E�qj�ş���~�'��Ov|�!�̷�4P���7E�
�T�'}�O]+�,OJ#��ƈ��o(d�z����oWb��<-��#R?n�0I~��Pcܿ"V(�$}j�1���?��:vxP����T��"g2"p�p���O���"
�u*�I�f�3G�b��M�;�^ԅ�G� Aj&o(RE�}^�x(n��d�J�j!,��H����'ݔ�̓�?�O�2ň�7q�t�`��6rny����;lO�0��'&���5E�"��t�����g���iH;fIՎ��m��L�@J��\����F�O(ʓ93��G/&��H�����	�����;qҪ��ɋ�T�����j�`��#�'���7>�	s��7U�h	Sq)�O�te+'����'+�� 0I�h:bq��5���'����X�J��@�AZVj�5F�$KO!���iD�I��i��6��O�����ɟ E���iu-iB��1L ��"'o��2�b���'�t$Lلڒ��(����G�z��n J�'�< ��e��G{\Fo��+7.8:���m�x4�3�'��k\a�tl#��OsB�'�靶m>�X��ʪ�T'Z�T�4��� .0zD�)�?���9]����C�+�L<�7 ('��@�SK�-|J��"��hlN2 M�K~���HlP�~&� ����:�5�!��4 �pt���?9�O�#����d��`ih8�B�ߠ.ܔ�Z�)	"~a�B�I�cf,�����SY\ �H6B��@�<�b�r���e�'t��		�P�P$�#��0��*hB.��g�B@т$���?����y2,�#K ����dh�X��3I'w�K�aD#2�8r�W�T�ttx��<lO�Ds�(A�}k��Ks��+hS*����'m����F�4�=��IxVxQ���.Ot�)�N�6�
% �e�O���1���'�4uk�n�=c����U�ɪ/��K�S�'�Iv�^�U�(@��OT�6j(���{�Eɟ-���͗uVV���=Yz"2�� ����Ψ0��OL-�&���'ve	O~����j�HPQßL�80�$�Zr�<�0��4<"q"`�P$JՊ5����X�35�y	+Ւz�z�0��(HX��ȓv�l�r!�²2�p��
px|�?q��)z��%�X�EDG�{���aND%v��p�r)͸��'1e9��i^x��O
"p��c���7��؎yҭM�D����}&�<2G��c���p�^��ՠ-D�c3ᄊFN]H]+sl�I���/�x���OmHP &T�T ���9x��J
�'uX욗����iB��Ãv�dk���N�$b/�ɏ].�:�Gp^v4��'�G5��IU��Ȓ���  �   s   Ĵ���	��Z��4��B��8�d�@}"�ײK*<ac�ʄ��I&`�r@x�en�x�m���S�b�'LL� ��H+֬<p�4|]��es�a��	D�F�Aal]�´BwJ.��A���+ww�"<��qӔ��ķbY�-Pt��5�:�+�W���fd�?|gЕ�p�/?�bŗ47�C{}�A��D\��1H�)l:&� T	�L��Lq��ŸW� �
F@��<��̌�/��cE�OZ�7r�� *q
��l�ҩ��_�p7 �N5\Z�^����@ǈC6��0k�<���&��z��\MK�,�y�����X.&( �#�>��I�3���p�Cn~r��u,�mZ��D�_�`X��׶{��(�u�ֹ���O��:��$H?{���&̕�:���G�����Dxb�Uc�'O�E�'����� �6��W���J� ��H���7��2qOXe)�a�

^Q���ey��Ѱi:6�GxbJy�'SL#g����t��F�9B$z��D.���'^$mDx"�K[~��2��0"Dj��%� �1!F���d)�O��ي��[�ƹS�\4,�&0� ]�{/(�Gx���Z�'�@�	1y7�I��
�o�@8&!�x��c��;��I�w8�'?`
`L�5��8x2!� ���'�TFx��}�ɝ�?���0B� E��`Co����Z�z�� �F������C\a���a�P�x���8_!��&ήu�*t��^�:m �Ő�@wh]K5� o���'c�M����T�'Wڵ�O��0I�9[2H��g�$gب��2q,d�A2��&$�`�"iۑ����$L	 F6����&D�`H��   ��pyX�Lwݡ���<I�ꟊd@Nq礍7WF�h6(�
&B|
&D�O�d9Gb�byf�O��s�Ĝ�*0���O,�D��_�D�a����S�@�����9U����O˓R���C�%��?y��?���{��ed5qV��sGH�FH2Յ�P~ǯ>1��~�K����*Ϻ]���,�n݃7���iȬE2�.B	98�{s�őim�i����uI��ON���i��m�0[�ܳ�f)B�n��rk�
+\D�%��$�?)��I�
�t:���?�'�?����Ĕ�V�lQՠğe���B�_�Z��}�2F�0}L�d�O�l�,t$+?�WR�,���H��t���0v$��`Ȇ�!I�I�;�QC�ː�z�dr�P�!NQ�v'�i,j�cd7O��sW&k��!�   >    :IZ@-�nkZ��&C�'ll\�0Oz+��AI��e���X�'iD��  ������|+�i���?��   �	  �  �  ]"  5+   �pA���D���\�'ll\�0BLz+��A	��e�2b������Z���'����3Û�� 8��*� [��i6ȃ�_�հr�'*��F����1-SB�P�Џ�'\x�!���'|���/E�9^��c���2!�r�E�?Q���䓬?�����'w����I#��]`���fHߓ}�'�lq��h7T�	D�W<.��y�{�Ahwr��_�D����03����	�Nd@I�=��'�f�;����'m|�YO~r�E�b8���uCC�0�Ȇ
Ok�<��A�%���F톂?�ؼ�m�]��p�?ɕ��t�����%S>Mm�`x��Fd�<)��Nh�)��<hB�@ �M]`��L����^$6QB�AJ:u���h7�D�y8� ����	2k��<�@��?xeK��0!�a��U	��@E�[^̓7��A��+�3�$D
{�T4����Ju.�#U@�0P!��΁C��EP�j�T`�ER�1O$�=�|�eDCzllV<N-�Lc�.Bq�<Q��U�-�N ȤҝT�q��=�HO�ʧ?�O��:�d�@D��Uh�P���G�'5���;�	�h�v#|rF��3y��I&oPeqX{���b��X0s��K���贀[b�h��WNR��E���)D��3 /�>o�j�	sL�L���)7�#���<i3�-d(�$��N�W!\-�S�TG�<Ic�J�DB���`��<Mv-z7����4�OT�GzBE#�G�/�<�"gk H�i�$J�Up�R�㈋HR�%�	ğ���ퟜȴE_�_�.u�	�|:��i�h�� �h�����[����-����O. ��D�+_�M��RWhRV<���[� �L9�t�F,S���R3��3d��������I��'2�č	M񆜚��9*�B�x���/8��{��&��ޠ\ߔH�G$�sP�mR�^\qOv	���O ʓ(�)Y%d����C5��`�u��*�To�5C��tD�i#0ɓT�d�(c�T�N~�t���C�R���+He������_hX��� Z��'޾5!�������2m�yD����31P]�Iʟ0�'N3��Q�0؎�B��
]�te��'��'��O�\]i��۽o��-��h̄��V�dPd���	��Ĵ����| ��B�5��{�j�O�˓h
��&N@� �@�|�I���U��!#9�������G���E�YQ��K &n""��Yܧ��b���%��C��8*�q%��R��2�S�'B*�蒑�ZLXs��ѽ[�}�I	jUf���O�|��q�'��d�`m����(��
C�nX����;c_x�P�(�6+"���"�ZC�'��)(Wz�Oe�0m:X(����ݡC��C���6�p�������-Z��R����������I%]R*��Ԭ�=''P}�k�6c�,eZC����Y���>O���
G�޿d��z��0�V�>��I-��H��-K�����Y%Q�t���(E�Gq(}�/��V%r���A�-�ҙϻ��) q	�X��H�o�np쉋�y�,���O��2��O�	�O����OF�wӊ��W���>���@:4U�����L�'`��� f7���(�"���)����?q�?Ov��0>O�A束d�P�c���Oڵ��Q�
]�b�ƃev���Aɨyf��1�1��!b� 9
!�4}B��)
<��"�3ج��N�)X�(C
�'M��{eេ-a8�H�b���pD
v�G��xa_(4A3Ǩכm�5�$�|�X����<��~ҍB�?+XH*���i�zL������=1Ґ|R�ZD�e���[D��8�����'?�Q�E�|�/�3>��[�'��FfD9>�6yږeڼj����F+d�d�O�,H�Ł�lMr���O4i���1|��9O�6mR>J��Z�(ms���dI"j8ay� �b��c��	t����� �j��7Dԟ[��DR�� �n��DȨw�b�'b�7�eӈ��� B0����%E6F�¥�a�Xhy��'��O�);��)�4�$f�!DA��ȧ��:��O>Gz����CB
�F��р�1�9��i߶��<Y1/�vIp����?9(��
S�z����$z�*�U睮� ��t����	y �B i��B�
�R�$5�l��I�j� a�Ҋ��vM�`�Ӂ�qQ>O<�ȥa�=���@+X:{;�]�Dh��U�O��u����P]x��BU�y@�L<᠁��H�I��Mk�����d�뎎�.6ʈx5��k��j��&L�qOl�$0,Or�2`AC�TV�7�dS�D�g�]i�'H��@��n�oj�I1y��H�IA1 ���
�^��ǈ��<	��?���H�N�.�+���?	��?���,� �8q��;�Q�g�U@QA�ꊗ��'�r�U��P"�E{R��?��1��ś{�n��u��:>� �kP�>ѕ�O\���'o@=xT	ҥBKAɦ!֋x��`k��O����On���l�Oq����+ք�v*�)2�˚Yr��ڧ`߽�xB)�>B� ;pc QA��{���?�5O�ͻF�Iĺcf�'����Ty�����ݥ"64kC΂�	�9�Vƛ�l�mZ��?��?q� �#U�Q:�����bմve䥡��Y
Y:f%��H�^�� ��_�L��$�<P�%��40��8�Mfܕ�mp�K"��U�`��B��Y��l���@�'0L���j����'447Ŧ��Ty��'p�OD9�P���\��(/ڼ9��'޸�On]� ͛�.�*����K4���Ӣ�DǻzQ�<!�������MC�e Q�2���J��]x�0��!u�'mx�B��9�R1��)��5@\�:,O��ab��:;��Ty"��/i�8���'%��8�C�-16�'�:�-�A���	4� ��S�5�d��	⟸�	����b�/!�n�ℎ�T+�!��-����Ob��?Iy�e�*))�Е��O`��AP�=�I3�HO��Si�uy�@�y��u�B&ۉ]A���ԍן��'������W��'��	|��AmZ"'g���V�C�uf�%���|�L����?�WC��R�84ctn�{~��O�~����P��?��h�2'����U: 4�'��N≿i��ic�J�$��}�R�,��')�C���E�*�P��CbA�-�'V�-{���?��i{"�~z�AiݱXaA�I�V�y h�,p�4��N%���`��I9�4��pd%����ίbfLQDzbҟ��ɵ����$����P&I��{bL$��x��޶y�$��?���':���ƃ�?���?��K@<������i��Ɂ>��K��<r�F]�Oh���c	P�vE���$K�]<�
���'I�#��Q��H��d,}r	V�Gq�c?O@�k'���4,��	BH��!QB����I򟜈�)�>��Ms�I�&>�(���'l�}���3�!��5���a�+a�>���m���o}�@�4�u���O��""=��+\$R-�E#��A�;�R]�DV9���V�g����f�v��M¦aSkrbU�"h��B�I�.���)�	DmQ�H��vܶB�60[y"��
&�Bx��51���ƓM�n��hI�g�z<@VS�<��	��;�}آ�)
ލ H�m�?A��3���K�jn2�kP`S��`����ZD��O�=�AHh1O
	`�������_��!bo�2 � (�T�V.�ybA��Q��h�GLh���ʜ�0=��"��9Xt4 �(ݽ5s*ɪ��,�y#U!8g
<٢��+���[���'S^"=�O/>5)�ɱCx���\,bE� 5�B�d�#w�$��@D��'��&z <c&	��
�i�%���K-1Oуa�X����t�r!��M&v��G�?q��]�ȓe1:�1P�Y�9P���H��K�jD�<a����×*�ISV��F���8WD!򤌅
,�U�M xzl�B�X�&�"=�(��(�?����?S��!�q-��3=b��5$�ן������'�I*��i�(P.MK�*��3q¹�hE.})����璪u�����?������,P<H�J
3�y�I�,��@�M�~:�Ъ�����O���\߰�)6��d@�:�ٟO�!�$��3T��M'g�l!�p�&<F�>9t鉷��p�����ɒ�����Ȅ4;ԕ����#��O̓

�} g�_�	�YC��.F���B�ˍ� )B�2J���!�jȐ:0\�Q��M�4C�I�L[A�FN�eQ>e�P艮y�Pm�ƓEΦx0"��u�\
QNn�h���~O�d��>w��!���K�O���?�U�3M�b�U���r1j�'N=�8)K�7d)�O�DR�R�(D1O�Ȣ���Ԅ
�Q�p���n��!������@��y����q?]#�`��B�Qt-ѫ�0=ɍ���8E1H�ʔ�G9�� �C��,�y"ָPʦ���M��T8��cC��'"�"=�O
��x�ᔕz�]	׭U,c~)hQ�6ғir����$�Lx��O˧^:��0���2��9a�1O�E{��ĸ��S�? ��R�E�u7(1��Ccɔ p"O���׀F�M��1QR�6����3�Ş���'��`n��%�B9M.�ȓ*�H�'l�$-Nf��֢��u��@���|�����OL�ʒ�ϞKw��IǨSR���SF c�T�T�%�'����dۺ^�LضoGD�=�7�_4K֢\��	y�*���J[(-h�Pa��<U�C�ɱQ)���れ&L���)��L-�"<��^DL��/=�Z\���W�Vf1��Hj��"���t�4��e˓p�FE��8��$�s�'R�O Pұ-K�
� ����c+"����O�=b(���1O&��g+��/��'���Ib̠z����)��;WJ%�'�n8�A�ACd4  W�.,��)�'��0�' @����Z��E�.K�E�O��L!xd���s/�7t1y�'"��O��x�mēV���k�P(ku�$N�'�FԐ���OVk�(��d��i���d���9��>�)h����<q m�q�ӎ|�Bx�������97�E�s�4D��K��؉IXh�w�I�PX�d��2LOV�`����gGS��T.,D������t��NL��S2!+��'�HO�S�yCv���aلe�:Ղ��5��h��$�;^Ď �<��&S�?��W��=�0�'�(3j�R��v�q�����%�3�䟹K��I��N&��M��I!�$ŊUJ��³�F&"&5iы��X�1O�=�|j���57/�i�цM���G��o�<Qw���f Yo�  t.��q.�HO��'��O,\B�,�2/�Xl� J@�P*����'���`:�	8��"|����F���JJ�xLZ @�I�?�N�j4�LO���1n./��d��D��C�/&D�� ���hk����D�\�H7f1���<1�$2�qڲ��e�2�XC��B�<���	���p�+E�;s�5З�����O@Dz��?���p����3&�=g��l�2������:-]ĸ���#�(�'�|��/q���5�A248�#��!�ybL�#W�̓p#�	&�J9�V��y�nD?�Q���֎��(�B(�r����3S���G-��</�1�����2��{�j.���.UN�
T�;�\� î`~�Of�Dz�K���č�\�H��GDI�wj$`����,K��h�
�ö#N�\��m&?Q+���OsTT�4)�:��Tr�%1D�({״`� ń)ѐ�[!-�72:��$-�	��]�G�?GT}z�G[ rN�B䉫w���q�ț19Ri��
�㟘���?[�(�� _$�'`�$6��2�B�HO�ġc'�o�G`��2,ժ����Gm�I�b���n��<��`�n��>�O>%06E֪R��D�#L6N��R"O2�
�&�-��8�aP�^����D?�Ş .\�Į�z"�5Ha-�4���D�ӌ�L��Q�^�+��Z��ĥ|BB����"y6��@eZ��̱T�ݨ1���6q�Xb���A@2§��٣G#_�P�����&���3�
z����	-w�`Ͳp��=jwV�K-�/Y�B䉎q�T(Z��¤T4�D��id"<��I���R��f�R�� �n��E�`лW�T�I�@@�ǅ?!���I���DBo�'���On}p�c�qyS�j���4�O��j4'D�1O���4{��O,�+� >�8U3Ն�
<�z��P"O���$�@}���AF
�6M`�"O���� a=бʴ���M��84����f[�(a�u��J�f	<9b!�7|O�y'��K�U�z���s�ԵS[8TPD8�	g�'�U���O:��⃈�\sd��� �/y�$ȩ��>Y�e��_��A�<�V�Qn� (f&��G�2L4����U�%�DC�)� ���T��aT� �A\7~��a ��'��O~�!�CD#l�P�!"R��(�Q"O�aP��C%b���T����DHS���i�@��2ჶC�t��tӻV�
�Fz�G��}�rb��pSh���ۤg��SJa(v�Ԡ' �m��3�� g��l����|R�A���4`�H${����Kǻ�y�c�p=)aԾ{�<��fߕ��'�ўb>��eI��|	��A�],��p���,D��൬G�[WJ�{s(�;(d�D��Zi�'V���'}��z�O�7o"���A��'|^@C��~I���2x~>�Y���A��3du }QR�@�'9��0�2�O�,{ulIm�Hi�Ն�b�ܤ�"O,aä�M��́���:Wn�����	nx��aa��-;�X����*���QA?D��Y�j��o~��!�ɒ 雷��O�`�'Δ#=yR�|rݾ,�� �B�9`?x���(+�~bL0� �y�#�O4�J>1f͛�R��ҡ;�V�!5J�1'_&B�	�g%��3cE��#B$�Ƞ��C�'ʌ��NM��*�nFR���I
�!2��ơZ䄈kL ��	
��n�"�X���|��Z5Jإ�F�?��鉚k%���mcr����NϘ���]�P$�|lڛH�1O`��D��d+ș&��Pqu�ǅS�2	C��#�y�
�-9)@�3�"�[�P�3�/���0=q�bm̾Q>�[ "��	uu�diɱ�y�)Z�[;r�{�A"�5� @���'"#=�O�.u뇦�pl�4�q����̐�퉾4"\҈y¤���B�%äf$�1����O-Z��wfU���'����s�F�g�	o���Ս� �0��M:zZB�A�2)Q��͔/;"̀��	�b��F{��4�ǔ	�<��:Hi8�
�y҇Z:�69`"d�d��8`�%�6���L�Ō㟴�R�W�r���%�	wP̅a��O�uҰ��R̓oux�E��NvH����ï ���(�J�b`
��dg��?&���x$����a�D�듣G@�<�f�/��uH�ϔ=(|�$#S�x�'��yrNU�\�r�2wm�2
ߨ������yb	"R	�U��ƨ���a'hW��?!�X��!����f�.���zq����(�JN����ɫ+G2�©.�i��ơ>��Η8T�0�qїk�Xi�v��$�!�Ҥ�-i��8@�१�5a!���I�~\��Ǚ�L�f��i�q�C�ɔG��hB��تX��3tCT!>� ��D�]�	�"�"H�h�%L����(��d���`���Id���!~��E9a��6
�KwHE� �On葐��*Ę'�nhK~ZuI��ı��X�5Zn=84�S�<��߲2-+�D�:w��B/�i���?���5o�mчM7�ؐ�p�c�<iSl�Dtt��1d����`��"���'Y��(g�Bk�*����J������0E�4d�<��>�r%ASqz8yd��?|_+�8;�tb���&g�8{\q��'�~�a��	�$��qC��D�9�+T[�<"�ͤ|����`� 6c�dT^��hO1���S��(sQ��CE��l� #*O ��@������ïHy���	M���'�ɯ>a2� ���e��ŉ�f�5ܒ�$�u�<�.#���Ȓo�8���@�W�,��Azw-C�,y������Xr�P2/T�o�@{"��-X$B�ɺ-$����&R8A�`��`�	>18#<�ϓ
s(��I�)�̉� Ō�q���ȓ�6�x"��(#i�8 ���'����ɨ���Y�'1O` E�2c|͡&��k�P��3�O���ъn`1On�;F���'�$'����� %o��(�w�"D�H�񄞵T��6I6���p��!D�� 2�I�p���1�;�Ua�/#4���Gƙ6)�ny#@,%P.���� |O�P$����A�c�0���{|T�Ã�J��uw�N�?I�G�EwVB��W�AP�EDl��c���`�%��!D+�c�!ߘa� Ǥ(�!�Y�a��ICWJ�^�X2Q��8-az"�䎦n ��Ş#9n�L�5�ٻ!��WL*`Ja�U�h����w��O��Dzʟ�90!�ێz��lr��\�o���P�7��uA�DY���\$���K5n���'L��1O���/L�Ӹ��P�(�gAV�K3eB&��}�ȓ	��!���&C.|5ÈN-V��<�����)������ b�T4�!�d�%��42'���d���2��?5�#=�-�Du�?�0hM��[S��6��C��\�9��`���?Y�!V}��iR�'�"U�P��V4�� ��j�;���*)b�.@J���>Y���7gw��t�;�L<���*��Ը�@�1N��q��=0TLɀjU}�#�?a�b?O�A&���TFA�l��_���35�՟��'�L%!��|b��W�\����'��"�e	@"u�!��I4}56���o�_��%�wɑzXRkc�t
r(��?A����D˵L����/�t �s	G�Jݴ  ����M���?)���$٨E����d>Q��c��6�F��ԡ4���S�.J�����4py��+��rx��`c
v	�eP�$�#]�d)��O�s�-��x���[Kx�0ʝ.�
��߾t�~���C�1m!����O��=q�}���wW�������oa�!8�����=��|2`	�-��H��L�e����&ٶ��'�iq��'S�I�0��د�06-���u�'e@��h�#L#(Ò���dyҢM�p�b1�Ρ�Q���1Cu8��ǫt[���"����Q��o�@6���p<�v��)4( � ː)x�"�a�Ñ��|zO�w�Ș9�Gϖ>z����4�y�'��ɒG���  �Z�U�^ћ��˳Y���І�ɬ;�D��r��g'h��6�
�cX�T���T?!�!ʞ��%�`�9�e?E���Ify�*�/����C9��T>�Q�4�u�O�^,~��V�Ԅ�j�� 	8\�����Oh�Ҏ��N��#�hEbI��j� �	p��U�tCf(t�@��|��� ���ēvv�]���v� 5�WHE�(���i5��l�Zժ�/�-ˀ�9F�x"�_<�?��h��6�A�
�(���(q�ޭ��k�>m!򤎓^7�X@S�/�1p$+M�}��#=�O�.U��B��6�@���Tp�Xl��I-��agNߋ%����O���G����U��0��u}��H�Cֺ91�&���h�ǝ?E��P1�\/x�')i�����"uX���'}���D��]n\8��X����e��,�v H�����������A�p
@5J?f��4fX��hi`q�'��	1+j�4�H#=9��M�愫��[�OD��Q礐E�<QH޼c@�*u��>\�;hD����'�V,���O�,�$�>�f�Ђ`�*�$�&n>�P�a��mY��
u�bӤ���O��$�<�
�?1�O����!ǂ�2�������m"��Vl�"*��S0m�
O���Ʌ�P���t�����O;�T����z�$�(�EF؞���G?�����X��Ӷ$�4�d�O�=��}r ^3/�P!0��1|p��c�"��=ǟ|		�2�lH�������ƨ��'��iaD�'QqO�N�
n�d
��e��u3��P	����ȯ��'-��<9PQb�ӁI�q2V��YvN\1^2!vB�1A��Q2�"*`yRD��,	�x��d1��.*fDɐ"m44)9`��(w�~B�	ka\q2G�A��up�AúJv�hZ���?��FHU�6Pe�����2�R��F�r�'K��"E2�I:5K��¥8���da������	#�.c�����#S)q��'X��hu"�'j��
~֘1
�'?�U���Յ(�t�u䋢{�t�Èyr�)擩DY^M��A+Ei�	j�/\�5pB䉊r~@(��T~�9x��F�P'�Fz�X>���2�I�ܹQR.��k��7b۳w��d&�O��H@  �   |   Ĵ���	��Z�Gi�Y��8�d�@}"�ײK*<ac�ʄ��I&`�rLxRaoӶ�m�+�p�� � j�vzpfY2h
�Hش8W�f z�-�2���ǻ\���{�@��i�dA>R��#<�P�l�6!ȵe%"!j/XRD�my���i��P�Q��$�PhҬ��4D?��=�^)�V�C�aø�0�lc2pA���nt�
���  ��D� PF�cEǑ��?��O��	`�bT@��!����!(�|��boQ	JS@\t�_Ty�/&e�r�Q(�����4��  'EJ'O��uY���tq��E��W@ԃtg��$�g C�+������=?I7��Q��6��M~b��1>��i�-@WL%2����y���f�'�� Fx�c�=m̉�%
�:-x��*�Nd"<��	>�?�����2d�$c��ac)��%��y�O8HK��$���'h� 
5,�y�2�ۮ7��q*ش;�x"<�u�+K�y�`pYr�yQ��x�8,9�iE|�qK�#<�0�6?)W�\�ZFPz��>&�Bb�sy���W�'����?��쟳D�P$0��=K>�@q�ڲ&� "<��D&�4d���}O:UXDA�V��ta��^�g�1O2u���A&��I$| �� 50�u�R�W%����zyV"<yV�0��/k�0%�|,pi��R���a���"D�2�ЯB�Z��v��;h4=�á��,�$�������<F'��$G:-l0DCqJ�:�\���U71c剞
��dJ�%��Y��t���x�*�3H��X�d����e�ŗ6��)b�*�(OP�ډ�D
ng,�ye'\,p	��{�B��!�Ā�C� �  ���m�\&>���O�%��H`5GD�-8)
f�Y��M+��� �;�@��	ɟ�[7�<�O�H�i.a��-��DRNC�*ǴiB�'��	��"��L|���ʢ)�'=ȡ��F�l�#L�qy����h4�	ݟW�s�l%��Әwㆠ�'�N���PZ�+�_t%kٴ���͜>,�n����	�O��ɍoy"(B&c�H��p+�?!�2�������8���?�
	��?YH>��GM�ӳNe@��$�M !@��' H7͚1_�*	m�ݟ$�Iȟ�S���$)�y"ĩA�����B�
	a��
/��7�Ve(��<���741�
���T( �T�YrH^�YBE�"Y*�n�ȟ4�	˟ AT)L���D]�U.�'}�<�4/   >    :IZ@-�nkZ��&C�'ll\�0Oz+��AI��e���X�'iD��  ���SĻi�b�G�@���<   �	  a  .  �   �)   �pA���d���\�'ll\�0BLz+��A	��e�2b��+!��/f�<�'��X���׾Y��W#,�ҩ�(+A>��'�UzÍހ
�Ҁ�����L����������'���cb`����p2#S��ph4ʉ<�?������?1����'Bq�')P���vǑ�$�͛ߓk~�'2�����t"q)ՆY?�8��{2C��I������P��O5Hu�u�W CR�`��%bg��O��sJ��H��b��SP� �i�?F4���9-0���E��*�!�dJ�k*vX�����{���fG�C�az"�$�'*��!�喵rj���C��!�dG1>5bW �$;{�!�&�Ϛ9��O�EzʟB8q��WX�Qk�L��-��8�h��H���	:����N�Hs��z��E �dDCʚ\�1OD�CʞԸ��@���fˀV��(����y�l��)b�����C���Q`[�!@��<y����.�Ќ����	؜Av�W�w!���~1�i0��dDӷ�����=�O��O8���	�2i��C4!ټFN4%��7Oȱ�d	 �	M�Q>�д�	�~���;�7Ѥ	�
-6�P��'ҬE�I�#2�r�r��ׁ�nD�'�qs�$X!k�)��������:<O1��іU��a�eG�!"�ɊQ"O*݊T͏:w弌��E� f @��'�8�,��`YM>�pD�a�Ƀ" �
-i1�#
5`��7�<pb�'�R�'X�u ON[R�'4� ��-�u����E�,L=�a�Z"
��X��V1�p>9�D��p2�J ȭK�ք�!HO�oj�P��)=�Rl�h�$/�,ԅ�	0.EP(��N��O��b���y�*`�B��O&�$��]��Dy��'��OP��炝N����ώ�n8�8�A�>a����}�	�?>б�E���2Gl(���K>Y0m�/��_�H�� \�ig@m����M��rQ��ҕ	A$��S�>���q�"		O��"���Y��O�){�,H,n�R�z��U��˓y��	���/��8�`xs�6{(�c�.˴9ay⦎��?9����$M.f"P�C��Q�a��)qgm��94�d�Oh�(�)���D/L�`Ơ�1��)iq���8⟐��T?ف�,�ʸ)[d�_����S���a2��	ry��)Ȏ�ɴ�Y���OK�y�;d�t��d`�k��`� Q��IN�H�`�I�t�ɏ�T�xbb�zPHq�!L����"��-�Gx��D��>Hy^dJPGޥm�D��F���J�B���ߟ�&?�&>���#�qp�͙�<A���-0ʓ°<1uM�OPت�::�p�����HO���k�v�tv(�&[Ȓ�*ȑZ8�1�ǽ`�����?��)�jtf�?9���?�`�ꑪ��K�x\��w�2@M��R�ϋ
)^0`��b\5Mg�j�f2f����g|��#}��A�fOL�┧�F�7���k�4b�X)Fu�3)Zq(-ipB/擎CLV%�wJxR!J�.B�ա�.:<^�P�$�m�I����P����Sӟ���������钢�	?�� ;5��9T��,1������O�������i ��4��-z�J"I��C���~�T:ǃw���3*?����@�O!�=�+5%��]�(�m+B�#M�F�(U�!�<���*&�fE�B�Ĉ8m���`� �TĆ�0��/KY�D�EO9����{�zfρ7dQ�l��2gk!�d��Q�
4L��FX�ZA�2���';���L_�0Xr�h&�,z�Y��{�"�dW�0j��c��7�*l`)�]�qO�͈��!��ײYi��(�'ڛ��ʻ*��� 3+ܱ6dp)Pw�M![���d�O6�D��0���$�O��	@mߨ0ej�9O06��[V��A&T�� ���E�ayGO�Ͱ]9��������	b{���4nL�GT=ԣ_0t���D�T$��'�6�x���(ͽV��<r!�Z3,�"\�gGAy��'��O�9��cy���!_2v��� ���W��xD{�O����ƌ8A�LȀ��Nr�fh*��"Y�lp�&ʔ�M{���?�̟��i�J�q��2[�x�#N�JIZ��r
�O���I�h^��������|�R		�XUL�$P��f8A�|�x!���b�'��usS�>% �#0P�[��`�ٳ��',	|�D�X+ibXrGb /L�'�̸�.�O��������B���u��T�[=���ff �CH��#s����']��'�n][��-a�fty�`�8��}0��?)`$��8�MKL<q'ț&'��Dє�p���He��i
�'lB�'{�,���M��?I����� �$��Ԇ��m��V;0��*gEÿȒ�'3����NDJt�F{�ʻ�#`K�.!+r�@��'�D 
��>���=*n���'�Rq;����i���A�`��T0r.�O���O��	���Oq����U3�����&i�.�b�#F5��x¢˯=��-i�&�1�8�f�B7�y�=O�� !��캓W�'d���
0�Ax�h׸{u$�����!T�`�"��5�v����?����	z��>�a�i� Y���#y��P`'������8�D���U-]�X�qgj�T�~0��CP�d��*I�dն9v�'KT,��)�䙱)3T%���ڂ}J��I��@f�j�Ŀ<�����'���C�۪:[8��3��!�"�Z
���)_v41�
ƨ@NL̩q�X>�<��=�ì�P�'� �R�g�%��Ǧ��R$Z.(/l��Miu@�Ⱥ�^,�	�<���PI.�����|j�U�si:A��<!rN�=2OJ�;@��9�갈g��aX���dJR�`R��&���4�g���	�>��d���QXش�M���3jr����,u;�v@����Iٟ��?��e��N'4�c�# HJ�(�
�K�'cў�)^�l f�Ux�Hu�HS^����ODʓO̕��	ȗ�?����i��Yl�
F_�E20�G�\E��gˆw�`0��?I��T�C@��p�	�J�4��'���IA�¦J8@ ϖ(�Ĥ�H<�f�t���O�(m����b��c�����5rH<֮Z՟��	ןt��p�AΌY��Eh�f��לU�x]�=y��߰<��`� D�:�k�B�`O�������hO�逸s��O�<�q�Q�.�^5k�3"��\�gK����O��F�M>@lZΟ4��럜�'C �чHO�[>za�դ�]D-����D��� @�S�M �N�=��&�����?�(��a��II���b�=���ē	C(��daOy���M�
�Də��'n��'��p*1�����i�$������R�i�,�sp̌TF�NH<����0Ub�=� �ϹV�$���<�'��{��f�=�������b�&�+d#$�H�í�7@�I���µ6�< H=�v�|[��	�s��2i��]+a�D?�y�O��U��K����w뾤����y�'�t�jX�s�0_������ C������Qs�c�.�r�aCO�+|�a|�|��54���R'U�U:2�Kw ��0?!`d��?!s-�H����&�*}�
�+tnMw�_�~㞬R��$��2e0dZ��]'b�p��g� �y�%_�q�l���LމE�x%�㇘�0=��"�!O"���KŬÀǠ�yRIQSg X���4�@K�Ō��O��=�O��@�R L�P��+�/������PzqO��Ӧ\� ��hR�F
���ɍ�2e���=a��P,|���'M@���a]C�R���lW %R|��'ar�l�+u�lyD����y��)�F�.49fB!O� Is���w�B��18���b��)�Ψ��KՁ�,F{ʟ��|�I�f�p!GAJ��N���鰟�p k4�I6iQ>7��$t_� �M�!E���N"�Lj�%"�Oi@v�I�g�Z\�6d�"�n{@"Ob!BnU�*t�Ճ��6U1��tx�x�e�@
0�uB��Rx���&$3D��Q ��7�*�)t��1 PEqP)u�L�'y�{��\L?��FP<^���K�9���v��88��ɑs��'���6�E�g���&X�T:"�@	�'fq�e_j���g��W.rl��'���Ã�pU�e�w��DA6@��Oֈ�GM�����VG��y���9�'k�']`�`ផ`���Y'�$=��K	��=�����Xܜ�I�#���p��d�Mi`*b��j��.��\J"x�ወ�e�����ϭ7�2�ȓ6`P e�ʠZ
�e� >'�
Y��	����bX�n��M�3H��3�\T��&����2�����O�k� Ex��)�T�Z<�Z�S�eX�"n�C���Q�'*R(;�{R՟�y��N�"}v�'C�@̞���2�	2f�)щ�L<� ��H�-�rǒ`e*�IP"OT�YϏ�f��	Ǡߍ+r��"O�E�b�Ugb� �NN?����"O�U��Z�_sVac(�'_\��X "O�\ٔb��,�~�'���Zw8���OR�� �)�'OH����5C��|Y'�^�2[�I�ȓ4b�Ԫf�5F�X�I�2	61�ȓ1� ����C&�8��3u⠅ȓ|BE��e�2	ef��l��yn܄ȓ=�h$��u4.P@�g*n���ȓD��[�3Br��v�թKw`�O���'������Rp J����Hi����'/.p#�7�%q��&s�Թ��Y�JyAa��>�
X+��E5BGZ��k�
�0 聉J��2�`��N�M��/�=�塇�D��q��.X�@���	�/�B���;<�;dK�&4d����b0!��p|s*ı2����"M��L!!���m1HU�F��%�>M�t-��6!!��I;G� �i�	�K:�؁���Od!�Ğ8�jxЄ	E�Sz��ס��F�!�$ך]đt�?Sdl�#�K4$ Q�Pr'�#ڧ8Ú��#�@b��
�-:�Ň�Q�Z|)���(����.G�{_���qЎ���W���%@��-~N4�ȓ�p2@�7B�]����z���m��<2�4Q��`�q�h�ȓ]��A���cP��Mj�`�[�:�Dx����G	�X��h��[Q���VY!��݄\8d�0r�َIc0�k�B�+u!��z����"J�!1z4*p!�!�G����J�nv�H�c�N$t!��R��m��̕<3��xv�S�$B�>)�P���UIX@��&��Kߪ�'mN}y
ߓ&Ύ]Y6l*C�,���3c�9D�`�S/Y(+R��Ү��?�J���$D��фm� lx���-ŶQ�V8b �4D���޼��
1B�f�L�P�$D�4r�l�O��{Pk��J<��"�O
}C'�'A���3Ɲ�T���J��:ɖ���'�IѤ�݂��UZehޗ�6"O|(q!��e(&����@��h�g"Op�Ң��_��pB1��0^�����"O�u�b%���$G�\~"4�"O*�)�B��J ���l��e�	 }�ޣ}�CG�	��0x��Yo�U)�.[l�<�EC=�h�x"(_uR���}�<I�ĦTN�(�慈'��xq�q�<Q�@N�]k(���O�j���Jo�<��,�<e��M��N�(U\���ׯ7�HO.˧Y�O�T�c`��Y�T1��!mDp��'%�a��:�	�K%Q>]��#Mq'�,�� �D�s4�ϛ>�Tup�<�Oڀ�F�U<\?�݃5ōU<s"OJ�`��7+-
%A�I��h,�2�IJx�����^98�
��E�NTP�C/7D��R��
�:�%�wM0I2��e�O�'��"=ѷ�|�j���N]sJ�#z~�y�^�~��p�*�W��YAb�O�a2aA��-��� v&��mx��a"O�(R�/�Y,�1p��ʊ7h�$��"O��`�HL��<��U��7e���`�.4��Y5aX�B��p(�BH���`�!|O��'���1 �.G�4A�F3[�x�c3�=��R�'R�L�!�O��a�i����7�0@/20���ε��'S��HM~���M�g�"�H�"Z
A�8�xHI�<� ��Q�`��[�"�q��C.(*lY�'��O,|��I:g`\f��&_(��R5"Oʤk��+.ȁ��SQt!Q�dXl���ə�-��<x�Q�v?�1����,u���=Yf���E�1O�삂�Oyz��2�^9v�bI'zfh�R���|hā��L>ɂ�J�S�F�*ֈ�8*��4���R�<�5�y���qA�-eiv�����51OV�=�|�K�g�БQ��׎"׮��Q��H�<ɷ��3>��@��͖4hm���HOʧ��O��b��Э
ݎ�Coe爍���'a!Q''�I�caQ>�u�4d%�l����(� �s�B��? &L@�)�O8���K�:Q��,�!�Rg,l�z�"O�؃l�^�x�8��/xorL�f�	_x���� p"�����Yl���s�$D� z3(�*��ۦ
�2�l��@o�O��'I&"=��|�FW�\.8m�G�݃q֔M��^�~rj|�&���D��.8ҒO��sCΝ Kȵ3�F�f�^���"O�S-�A^��)�%3&z��:�"O,dTHL�L����S�\�P
$�-4�L�Ed��Q�����[3q��`�-|O��&�D�QGƙ-ZLȆ��Q��y��⟤G{N>����%�ތ&�^3Ƒ�&��MW�O�`��y"�����pn���L�*�x��2lI�]��Մȓ=�v��F�����:����P
&q��c��/ٳ�)�@��2-	By��TԪ	Z�@FB��<ڰ�,�I�?!��)�s!6�\��j�&nO E��g��hO�]p�h�Y�$$���|L�i�I+���r##`��<I�R5#n�>�O���G̜wD�z��U`jm9�"Od��R�Ԭ4����4%O�Ѳ��$4�S�'��h��bR�B6HpTʒ<��A��8�E��鉨o��E�ue�AR�}0���|*��DA=Z��h��n�c��ŷ!RB>9�b����t�O��=ۖ��=� z!F��0�����kJ=�j�����x1�̇9�����/[�5�`�ȓR�C��3u:��GX6Y�|�ExR�'�Y�#�2�P�8�iG�a��̐�'�V0ȵjI�(T��xAjBFI۟�9�Ov�DzR�)�L�/���F�D�j�Z�c�'�8[T���Ħ�S1B*�I>
X�[`�=��N 7��I �"
�J$�I�A!�Mt������"b�
��UV!�d���츅a�5��,��J#qL&C�	+kn���G� ��܂��P/@���H�I=���Tm�D3��a�dV�2�H����\�d7�9���bw0x+`D�6u����ӹ3��'4�����'��P	H~2�����h�CΖ,*���N�R�<�̜�a.l�!��Ì]o2�
�,QV��`�?9ǧ�1�����)����|�$@�N�<T�D7D	�e�:Qj6���&�H�C`���'@
��` �K���v݄-
�I���
=����<�BT�?����;��x��͞ 1B<���V�tjl��>�3�	�'��|9�� �੘R"L�!�9y?�l���ah:���:q�1O0�=�|�@.��J[)#�ͫ	T̨v#Fa�<aH� �4+ ",3�]�!�ӂ�HO�˧<��O�(p�+�`~�*P/ǏRJ6H�OV���#�̓J웎�IKYh���a�'GzL���c��|NЉ��"\��˞ETѧGhň(ۆM+�y���A� �`a��kɌ�(��Q��O0��$L-1�`p�W�*y� k!��;]T!�I( �:6h�=5�Ȁ�+97�/�>���ɮ��*�0���7Cv��x��$$(P��&٘J$#d�ٞJԏ�d�	)��ҳN�4'�����BALB�I�r��IД�Y�g��<�$���XC�)� ���jP;����GW�&x��x/.4�����bN�mp�M��J��H؇d:|O|�'�  �� /<!�7��/T��awO8�	\��u7A��?)��\k�YAH�b�,ɋƪWi��b�tzF� ���$��؛���jm��_,m!�_�{��8�Т�1^�4a�fi�-azR���
O(� b׮S>Nh�@I�	 �!��O!;q��W5c&��%	R���OV�Ezʟ��#�u~� �u�z�M���8�ro=�0��$r��Ԣ��2eU��vtJ�C�I��1O���cO�ٸ��c��  #K���P	�&^��ȓ8����g�]�\S��X�.e�<i��󉂙uò	r��>+�D��%��+�!�$D�[@���&���� �F	_�`"=�(��8�?1�ǃ&b�L�rN˟H�Da7Ɠ%x>$���?y�Wlؘ$�i�r�'���'�ts3,��F�^Ū�`�rcR����߈7��|��,t}��زH��<���|��x"c�&��maF,����M�C��(ȵ`��V���d�`T���~&��e��r�e�gʞ� b�"�?��O �Y����t�ɿu-�ڗ�'>�ܹ� I� )�LB�	�gE\u�@ڱ|����5�*3�����<10@^��JD�')�ɧw���*0�D�5�l�K���j��}"'��'[@���'Yb�'���5��DI���$+��<삤�ׂQ�^�𩋬L��8"ΦL:5��n/�fL�㉬��M�E�Da��u[vh��"y4�z6��i����W�S���Z��'�����gR�5:`���Ԛ7zD#���<����hO�c��`Wc��G��vv�'+3|Ox�&���e�p�R8���^Ͼ=�mC�{����R�D�IC�(�V��ʦ��L�`^Td@���1� @�m]�?��$�q���	�?a�O������y�8i�P�`�H5����3fv0L㥆/w�t1�� {8���s�ZA��� `4̺���̌S���.���ѱ�c[I��x�o��<1�����ǭn�ބp�S�"r� &��?`~qOd���Ă}�^�#��Dts%O׾b��O�Ez����JV�>-eK�խ~Z�m
��ۉA�f�D�<�#Z�-&h����OU^��&�iF4U(�hU�L��G 	A݋�@�O���Np�i3��\*:��!�O�T��E��Q1�'iW
�GΘq�����Ȱ��'�X����V|����ƺǈ�ҌS%O�D�,k��8:�h\�Đx��þ�?)���h��7m��t�H�]-mz�4k�u�!�䄐u]8�{7S���f�'>-�"=��O �#�eT�/�H���<p9��b��7EtB�C"O[$f B���OZ�H�0&�j�)�O���g��aBH���I�rH�p� ��Tԭoh�S�#Ҭ��Q�I)y��a��b�"t�g�I7�\��(�
�~j�	�C�@i��7O���'���sG�)�3��5V'�Ѐ���E�h�#�n2kHh���A~2��?ͧ�HOn�ЄOJ�m�5�^�kU�La<!�$S#n!`�p�Ғ7|�5�fc�z""#`�Ђ�F/��?]a����$�Z�n=B��Z*s�2�A`�<C�2����oY\��IџL��̟h8�� �	R՟�ΧPUV�P׉w�0�A��V@�9p�
>�0!yr�~a{��21랊!>dZ �ܧB�!Y�(Ƨ$ծ���/lO�p���p�@p��[X�����	���'hў��>���C|z��G�J�'8��f��^���L>�r-��"wT5#@�L52UiQ�V�ef�����'Qʩ:DJ��`���!�5ӕeA�8|�ę>Q��K��V8�<�&��@�('���A�p�����#�@C�	�%����F3͜��MN����$-��?G.�I�$~!��;p�C�	�A����͇p���3�h	�h �x���?I�C�C��|�!,��d�$	`Q��HO$*�Y^�	��S�}涬q �	*c?X\��튳*����<f%H�*7��>�Ofh�U��0q�<u�!�8%)��pu"O�U#��C�h��|�c�������D#�S�'d,� a�c�+
	��W�0X��ȓ%�XC��B�c�|i���?��:���|ړ��=E&и�AŌ|䚴񧆃L��D'�Ofբ`@  �   |   Ĵ���	��Z4�G)Ď;B��8�d�@}"�ײK*<ac�ʄ��I&`�rLxRao�`�m�+I���P!��,M�
@j��T��A(�4[=�v�s�P��#)���t�($�&���Cś1�8��"48��#<�a��s�!د3u"x��+�]�<�(V�@QG.�~8x�ʰ#2?�3�*B�7�CL}"�΂*�x2��\��	:��T)*u����!j)(�u��<�q@˪,�����O��S�'�T�rkWK	�+S�#K�H�� %v�!Q����ֶ3
������<q�+�G� R��N\|���S�5��ȣ�I;1s�y�'~�� Ӆ��LLƵI�O<��d���MkW��@!��ϟ~��Hʻ/F��wCe� �g� @�\��f��J'���h�c���O�����p��O������]C -J� ��>A��%�>(��<0��A�m S��.[�B�b�dn�<{��$���O�e���Kݩ�J�>)� �U�M�m�O�T���������sx�]�a�I%JE��y��l�I�&j�$K'�$�n*���)�|�(�A��M.t3�������O.0K��j�쌂b-�Iv�
F�F�_�@�<�A'9">O�QȖEM�􉋧n|����Ov!���®��n���`'"K�NWv��6K����G'<+HY+se؃mJ���J�.9d���B��0��=��� Q��Ş�Vt^,H�U����d�hamI"��I�'C��R㩅���'n�)2�aJ≭u�v(�B��Y�\퓥͊<?h�"�o:\�<�#:�@\���
a�$�4lP�1���^n�   @�?�I�{��!�P�+^`�i��C�$I��C䉻w��=�GT�}Ӽm���!:Ҿ#?9��i�%3�m�6�� ;X�
⧅�U�!�����1¨��Z9����e�_�!�DD;j�:h�v�(	� ��G�B�!�D�VVHIx�B>"��b%�;N\!��*~�.ň��ªr�\P�C�OO!�dV(���zE�T &��(C��j!�ć�X!������00���bȥq�!�d�TH�| �D�
)��9���-�!�5G@���7�۽�0��$�A��!�ĝ��u�@B�a���[ĪC�1�!���|˦�A3F��&�T�V�F�!򤀙,�yY�-�2^\>��Q�8�!���P������L�ITʠ!$��
�!��	,ږ�s�m�x��1���/�!�   >    :IZ@-�nkZ��&C�'ll\�0Oz+��AI��e���X�'iD��  ��ʠ�Ц�8G!�d�*A�   �	  �  (  �!  �*   �pA���D���\�'ll\�0BLz+�@  @��e�2b�0��������) �ٺTm�'�t<yÚ�|�0�{w)��[����I"n�l쫢�_(c�~}K��wǶM�I˥:�8E��ɤ;��et�->�bę��vNr8v&�O��%���O���'��&S^ AEe���:&-	4�����r�I�W�^����8�l����$�@�4�g�̟x�=��f!���1�Be-�-V�a`�JjS��>1��F9 -�<��E�]�q���%�� ��Ƥ�C�I�6�����h\F9�$$I =�����1�I�)T�|8E�[B����[R�C��<%}Du۔��+OgQæ��'��詈��?��+�:K����$h�(2�-#@�YA�'�.qV!-�ɲ��IY �@W�A0@;f�R�l@l�pb�H���\�Yq��'|�XG�\#�(��Φ 4�m��'+����߅SƸ�d�>x�yH�y��)��'Q~D
R�(	 ��0+��0!�C�I�J�J8�'l]3�Z*�-қ#Z�#=�.���?Y��G�!5�] #i�+��d�$��ٟ�����Ϙ'(�X��	���%�uN�I��a��)�f�0V�[�#����U�،x���U
��fD�y"��a'����gX��ؘö[ �O���D�&l�؈��˻C�n4��L��A�!�G�vr�d0V%�,S?��zЀ3�r�>1�����D��I
�oͬQ�ZʒB���I�+\L:Ś �'B�'��㘬)��+��'��KV�c��b�K�8�	vm?N��q�JA�1�f���$M�ѰbeI�_�`���#��_�:JGf�;9Z�bv+K3;�բ�/�z�����������P&�3���b�A�$�����Odoԟ(�'�b�d[�h���2*Y�7� e*�k.-铤�On�%�hÅ��u��)��s5�-�vH����"�-��i>�	�yH�dk����7S�����WN���)2J �7�9�7�Z���/n�T)aØ����(@fh�i�P^�����D���<�b2�X�O���V�ˢԢ�ӯ{%F�IS�'
�=1���?٪O��G�� ��+����,� Z�O�iӆ��;�)�%�P�h����hxh�_� S �h ��T?��`�DN4�i���C0`Dp��W vN`��^y���H\H8ajL��OJСϻʢ�����&���b/�L��u�O�H��#��:�Y���ğxB�X�(��!���7^>u��/��; x�Gx��$l�9�&��t�B+3�bu��_6��Wd��	��%?�&>qC��˷�v�Sčc`0��$�4�°<	G�ڲH�ȹӵN��}�i��m��HO�ӀY⟤�S�G�w���s�� "B��IK� >4��"���?���mޤ�5�ن�?���?i�_Ӑ� ���
dÃ�"�*Ԣ3)��!�
�)�M/�D�H!.5	��d*1ʘA�T�2}��
�1f��H�D> �f4	fAX!K
0 ��C��B1/k
�#q@$�ӂYyJ�Z�wϐ�O$ @(�#$�6W��J�LX����şt��J�̟��۟(��ɟ4�	Ѧ}���V���Š1��3;+d�0�%���OΔ���S(܀�;!oF��ɡ��
��v����)n�hZw�,?�R鴟��O��M��e�(2x��	K�~qn ���H7cr^�P!�6�I	<��Θe�DS�a˴L�ůT��R� �=]���y�O:�ʕ�}�Э�m��m��\�N�?�!�$��y%ހȂ�B@�XxBf��K��E��'h��䃷�v�:��Z�?�����a`9�{�!+��7�pt����k��@�i�1qO^-��-��΀};\)*�'��&�zX�������`�y"��D�O���G�]�0`��$�O��d�
���9O 6��1���Pg̥ja���T\"�ayR�x�&���X##���ə;?�qX3JM�?�ّ�t�r��DԚPr�'�n7�n�*Q�t���ޠ8��MV�Z�Lh��ty��'��O�4�D9R-�y;-�E"L�z��I�3A�O"EEz��6Ģ�OѰ�{R��Kf*uZΦ���jy�G�Y�p p��'��\>rܴ�M;�@��	�����lC�tg�<�7�GP��'ݐ�1D&��svީ�O���BM�8br�',���WD�EEb����Bx��9I<ѕ�ն �.d�R%�'g�vц��C8z9'>���Ň�@݉��J�a`>%���#�d���'ή6m�O��OxT��Y�
�����F�����#,����=1��˰<ٖ#A�Q5*|�����u˔��#���HO@���]��ش��`´S3�AO���B�N�5��!� ̝�yB�'��Κ!`�l7��O���O��S�? D��F:C�*�Aݬ�T�h�/���'D�8�1�MF{��W8vv��X���	*�h�JS���9�$�>�R�R%���'<rX���.�n ��"bk y��#�O^���O�$*��Oq���ͦ���
��a)����<���g�:��x"ķKX�����Μ�C���?a�8O�����[`�'m�I�$j4C&��{*ذ(H�N����a'��Sd�0���?a���?V^��y>��k�0(��1�c94�nQB�߾��bU8���ݕ�Ĺ�LH6
H��"ǌ�.��y����l���'��(�q�@�d9b���(V��"�ć�?1"�i2�6��O���?ш}RL��;f`�oԐ鰥�K5��=!�|��^�;Y��ID@;`8�Z4����'f�����D׶
�x���?�ݴ�$�2�!��k�C�5�݊��'�D@1G7�h���'��iɃ(���J`��򄇝'<ʔ��N��^��p��I�".�ayriК�qO�JW@L�Aagy���`�̰<	�d�՟��޴y)�6�i��Ec��ލOAZ!P�O+=�ҳ�<9������Ov��u��;B�Ly	`�3d�.�9�r�7�S�D��(2��}C�嗂PԚ�#�Eޭ]b^�����$ۑ���*Cf�O4��|W�i����ڹL>"��Ν;�
�q�� =	��$�O�� H�[�
,�>��Y�	�L�X��"�%O��y�<J8O̲��)���1�P=Hv�d뢩i�aրN(�O�A�e�'U��'���
��i��̻qX�`��|qO��D=,O�(⏔�A��	�� �<g�6�a6ғ��T�φ��'��P��;-���&��K��I���؉�~��'�r���l6-�O���ON��"M����+)^������Y^�U��(���9?�Xp����4Vў�����Z�P2�)��[���&�N�b>��Ob�� �U�g��(�xXy��D���Cff�U(������?A�gg4�Q�S�gy��i$�x�@@����(�SL��(B,$��9�-T;S4���F�/�u����O�͓!$��Dx��|x�Ic}҆�m�y�%��}�թFM��~b�}�r}!���ݮ@��}[K>�-B8l~��V�^�}(�YECy�<�a<"H ͑"AsN�I1@p�<�B ���D�vf��RS���a��(��xbi\9[�2�	d�����.#��=��y�� �LE�A�Ŭ��eE��'Yў��B��$�?���"0�9a��&����m�$�Rc�<:g�6���'t"2؛b�[��A�0(қ�!�ɫ$�jp�q���m�h�Iff�?�az��n
�9� �N-��P2`�]?W�!�D�O�p%�tᇶW�.����֣��O�\Gzʟ.t��>9��<������a4ړ]T�:u�d����J
]@���th��b��T�=o�1O����U$Ѹ��v�d;��¬����2��Y�(��g��Bv��� ~�@զ����l�<����d�1��Ŗ.����IVv!��f~�]J�'V�`*~�unь,#=a,�v}�?b�׍w8\�v�L	�l��cK���{'n���'�Δs���'O>��!h�4c�����)�F�bUp��ӣ5��b��N9�=PB���K��0*� �y­�G�x�F+�+UZ�9p�M��O���DȲN;$ܣ���i����˺�!�ĕ�qsP�rw�		_��� )ê%xbA�>����W�a�v-C�k8 �z�Æ''����C	�v���(OPтM>т̛���j�*�O6^lBg�S�<�Qc5��M�Ս�8Q4�"�N�Q�<!"惞k�i@�Q���9c�^���xrCF6 �.,��բL �A���J��=a��|re�4<h
=H&�D@���KW���'�ў�]=jP�d�=Fg�<�i��1b��6���O����y�M����+p�����P^����
�8��e��iqR��qo�Z|ꡲ�F��!�Y��IR��s\H��G'��q��H�K���ȓUⴥE�Rg?��*vb��I<��?Y��)Ҁ�)a����1HD�O��`1�ʉ�hO�4ؗ�\̓r���!��|� �! bD�K����T�i�<��Ho�\Ɏ�L>� У��ѽW�(���}(�{B"O���ꝑl�Tpؤ�ƺ��� �$9�Ş9� q#3�3rЉr@���b��-��{��X�g��1��r%P�c��8!��Ļ|j����F�8q���wɢ@ ��U��b��("Nfc���`��O�l���P��-Yte�t 8�ޖ5���$�"lLeZ��2H�рA�3V!�$;x(�j�U c�ΐ��,�EN�L�牁&����EǣRH����b;<��B��Q��0%�ګo�\��AR����I@}r�7ғ��'�����cH������	�GQN��'�6��%'bQ�����|rN]0JvX!Kޏ%}48� �,�yb � 7�xBPG���RN��y"`ŀoR�H���#�d�z�V-����F�d�v�b�`�_��4��c�	f�{��;���	$Z��A�Z�T��,�O|�=�� ��m�I�ca���`�F(\�HQ�D�sb��Q��X3�Ob+��W�X��GP�	zX=��'���P"�b���Tͅ� t�����'����Ǽn��B�I���p�H�'$���VÞ�B(4d�����2�2�&�S�4f\*Z��z`�Q)`����x�Q�X�V*&��/��D(��/#�aÃiI// �Щ��T�1O����ܪ����Z�PUI45lF�"�ɽ\Ƹ݅ȓ5H�$��KV H3�ȸejQ�y},��<���)�5<u[Ј�t�-�e(�*8O!�\D6l�ulW9f@����H,8�#=+�n|�?)#ʋ�y�T�zi���t������؛���Ș'T\�G���,&E��c�zr�W�� F��i�aB ���?I���`T&Y�A�̃'�(��#�|�<9�ɔ+j\$��V���z@�g�Cq�'��y��X�R��� Գ7:L����y�%�/.r4�5.�2AU�)(.���?Q�R��S��D0��%)�m��,ot,�Y��I^&�I��M�(Me�',lh'����Y�l����䬉7�,��`N/D�4@�熘B�L��Ǐv�����"D�D�Fvn���ͅz7
�1��Zh<��(�-D-�9bA�y"�[��P���0K>��Y�RH���v�X�t�`L�6�h��hO�Ϧ/!���=��1B��L�M1�=�	�1��''*P�<)DANB�SO}�0�$��#9��x�*�Vo�C�Ɋ4)����m5f�����B�Zw����$��"5)V�HI	�PT�L�f�ߞF�C�	�L$�p�C"c����1�z�賎��?���`[�x�>x���� u�	��ZP�'���#��!扔3��)���HE�F�y�b���M	��4b�<ˢ�vq��'����`M�K~��X�g�;�za8�'�Pl��n�W��`��L`�pz�yR�)�S6����Z>!*\�EG�O�\C�I�h�j|#�,Ȗr(�c$�%j���Ez�Z>����H!pp��LY�:T"�AT���?���8v71O�|���IڥV5t���M�9:+�j���&Y�E )��i��>^ΝbĭU�*�,�hq��yn��\���ǂ�*Md=�Ѝ�O2��$��UA&�`��h�D1�ĆH�!�<L�6��r �'BQJݠ��op�>��I��l`��j�DA�[��؂t'�wVD�����F S���'�TB��|����Q�u`�! tX3瓾�y�!S�T&nd#���5bT�G���yl٥+���Y1���D@Zq1�N�7��B�V
A#S�y� �Q�Ӻ/��{r.<��(��c�ˋ�j�� ��=��Oآ=�T!	��� Tj@��$-�b���'�e�<����~�S�r7<��f,�C��PB$
6 M�B�)� B<����))��G%�-:�e��'��O¤���'_/ %���R$�!�"O�-
b$݋��掌
<����K���	Q� �ڙ�7���	��	G�挣=i���	�1O�t�t�O�@U�2��.�QԎq��0���J>�@b��L>��)�+Z���#gMXAL�Ū7�WP�<�R
�����WBB�YJ��hO1���j��%Y`��5	��Bf���C"OT�{���s(�8#�I_��a�3ғ���a�C�0钀��""���������M¹puvc�����S��D�X7��v�]�7Gځ_JZ��MA������
W��|���ΐDêI�����}�!���D����*G�JZq����~��4��	+VB�t�faۺ��)�'�ʤ0^C�ɼ��ՐE��V'�5��gb����Qx}��#�x��'�FNN8(b�@�<c> k�'�6�Y�k�O�9#��"��G�-�d;児�F�<l�F��1�!�T��±a4("R����$�O	t�!�D�K�D�'��O��}�T(�+�hC�7���a�Z�Hi��a6wEX��d|�	�~լ���+H,�l�aeX,K5��D{R�Pep�:� aʰ`L0b����d��'��O�Y��yA��uP��I�#S�D-9fR�ąȓm�4x��,�������
ʞ����i��w�q!�&\������g���ȓL�)�R熞[��{��W+_�,�?I�)��gFl�d-!`$�n�d��S�9�hOh�a��G�B��M�ӿh&T��D7\ T ��a�%�q�<y�B�%��>�O�����-rR���6"זl���p�"OL���4N����⮈5I ��Q�<�ŞAx��!���nN�ik
L�=������`,0R��a�����CPH��$�|���DL81�g��,?H���g�Y��b�9Db���t�OU 	+ЎX�K�*����2e�Hr�� o�X|��3��็,�~%�Ă�R)9J,��(D%y`�Y.'
���' ���Gx"�'�X�pF����Is%)GL��z�'U"���Ȓ>�~t�$9.<����A7�	��HO�4$�(s���'����D��t�Ȁ��L��	ܴ0�n��<�f��0�"p$����+f8ԁ#5�������=D�|"�֬.b�;�L.��Ì:D�t;&Û�����Z d�;�Wh<�E��8/G�q��Dqބ��pHTr���N>Y��(\��K�	�t��vhr�+���̺����?���ɰ�������\��`TiFc���,p��ŲrK�O�\��v#�����g@[�´ ��'G ��0��6U�A�6D�#�j�1ӓ��'�JȂ �.��� !�G�4!c�'�F�YVCV��@�*цM�-�V����-=�S����h�8����&`"V;"�ژ�ў`���E��'�L�)�'?�D��T��)Ic�	Xd�NXTI �yB�ƯX*��}&��:B*�5+�zq����$d���)3D����؍u��ق������ 2�\���On�H ��E�`�І=TP�l0	�'� �
��W�9 lY:�� K60��%�Il��`8�I�P���fi��p��qq�	pB�D̻i(4�<����Q���@�X81{�I�=��|��OP�B���g�'f��*%%B�N2t��J��9#J9�'�84
��A!m�ԅy!O���j��'<O��)Q!��,I�b��.%�P��s"O�Pp�`�-R�x��#�J�"4��R�'	t�h����K>����%̤}����t�tx�Pu?	��A�h(�Y�<�����h��&���F�+�����ܖ7!�,
2&D�� m��oZ�S�	��S�h�p�6D�� :\�T���=H�5CM +LT4��I=4��Y����I�eJI)a{�3|O��'��A��	/m�܁�ǆ�!���;U�/��I��u����	.m��LYa�S�y7���.�:b�x����=��O��HC#�* ΒY�ψ�܈e��'D@a����4�{��۸t��)����'���T@��!�"V� ����'U�t�3kMM03�@Wo!�8��R�(�S�d��$7��`��J� 6#�P�S�X;dў���&R�Θ'b��k��i
�p##)T�� ���49^"ؐ�y�%�u^�5�}&��9�kŐ$2r�� ��i{��5D� )��Ixĉ��7:�vu�2k0��t���O�
4��)
	Fh����	]t�P�'y�0�`OJ�b K� J=P����It�d�5�I��xq��� W
=ڠhR7��!Pl�	֟䫇!�!�M����?����?���S��)��ϗ�&�S��߷R��Kv��h���>�V1[���XP����z�HIp�.݋2cRRh�5��L��a>\��'��@�j$�3�D�{���ʳ ?S�d%j�ƀ.a$X�	c~�b���?�'�HO�u�+ۆ*b�ਃ(�L��XF"O�����IGV���{�D��'?2�I�'�#<�Ӆ�?�O�d�D��hº���OO@�@E�0%��M� 9�ܴ�?I��?�O��� hEƟ�ϧe����C�� ���Y�� ��(�#�ҷR��9�m��U�!O��0�F�+7��jg�"�z��Ц�y������U�h�(c�1�p<Q���
yNrGM�<q+�cǋ;D���ş�E{R�䎷P>��Ya9��DD�{�&�$�~�2`3�Q,m�x�5���=qOB9AUk�O�ʓ)�x���|�۴|6���FcXms:������S�����'$2%�#hH���'�i�Wr�`U'��p.t�6��uX�-iS�T=0�<eං�gCʰ[�z�(0�w�A��H hUZ%�1��(�eg�ѪDA��]|�|X�m0O��A�'��X��r�h^�h���m��2����;�	~؞��wH-\��:abX7{M�d�i=�I�HO�� <g�8��h�&jC���j�QDtTC�m��,�'
б%ZJ���	Йx<7�3�prɰmu��#�\�.}��؟L[��N� .��AQ��/-���� bł�z�����K�}���,Z� L7��?7���*ă]^��(P�ӯ4��}����4.r4P#�q�OR�,��'[�>�mZ�r_����E,
�MH��S8ZXB�I�t�ZL#p$N0s���c�,N%uhd|Ez�џ��2T����|�d�a���'23HUY��!<�R1�w���Y�Y��ş<`�������������<4H��)DDT!��R��愑�L	LPQC�qy��	��F!�m�w��."D��ēdR22���$����e%��؈��I)vj�A��Oҭ��V�g��m#Q@��8B ����m	�+�T�@�����w�Oˑ�RW�P*h7.���
.q�ntP��7D�k0cſNb2в%�}��Y(�O<͓$�l0Ex��0�2S����Y�4z@jRKE�<P��;x��d�W����?Q��?��x�
@aRf!�?�O�6��QD�'�Z�CbQ�)FB(���+*(@��������D��}BE��>Nn�t�f-L�z~����S<DKFh���_؞l��MI�$i��	�˔"3���L�(�����O$�=��}r͆���P`�̒��<J4g���=��|�B F�,Òe$l씸6��.��'��	Br�'qO�-�Ad��?�"�K�U��E��fM^�q#�#}r�[�m�|�x�y�E���'dW���'(�h���ۺ0 ��ȓ��]�����K��u��\F*%���_������C	@H#P�t�&|�ȓ/9�} W%��N\x��y[���?I �)j2�F#f��5�cZ+߰Q�1T!N���|J�L���'� iB��8���s��4�ԭɥC��2s0�وy��]�Us8��}&����ņBX�I�+ʲ}zz�JB�/D�,	C���O�vA����W���7� �	X���OO��s�� 3]<*�If�
3Y�}��'�4��	S�>R��¦�D�(���X�d`=�ɢ/����B��ly�"�� >C��IZ��4�ը�  �   {   Ĵ���	��Z�G	�;C��8�d�@}"�ײK*<ac�ʄ��I&`�rLxRao�2�m�+|�a���!t��v�xߴ�&�h�0���	.�v� s��^E��⧛n8��z�8#ϼ"<�ufӐQ�H��5Sn5��+RԶ|CZ��arA�	�DP���.?�R�Q��6-e}� |!�"ˋ/ �`����$@�4�P�W�f����PJ �<ǈ;d�%sV��Op�ӗ~�@H�C��8L�MU���:!!�::�TxSU�,#�Ra�"�g�<E��V4��3���=uV��J	�|D!�F�Q. ]Z�'�����v�B�9?Q�U�3��7�Em~�d�62��DCmφy,�E@��X!�yBC�K�'�htFxBbS!�XMs0�\�MB��HΒ(�j#<��+F�\�xd���c���>�<�a �L�r�O�큍��Z0¸'����ңu���C��4b���޴#�#<ipd=�p�3�!خh�f<B#C��-4�-�v�L�D"<Y��>?"�M2[�PDAU/��CC�Q���Ly�
�B�'�\]�?�� 
:��� E�1�\<��cׇAp�#<7�1�"���d<|$-�p�hR��� ·5b1OP�p����ē!�� �'�&a�-��e|���~#<� *�$1#�,� �hq���.��PV Hq���3��7���pX7&���W!K�c7�ax��'f~6��u��h!��'d�ʰjX���8rő�b�d�,O������Kr1O�ivL*��8�C�Kؑ(LVt!�[�Dݬ��P�T9x�Fyb��W�'�D��rJG�w-�qPu�_uxH
�'�:aI@ ��Z�R��@"н���G�?�*O��O?��S�?f�E�S
A�
���cZ�<9��c�r9�5f�":�@  O�<��)@�v��H־4����N�<�0��I �	��H�%���H�<�rL�4E �sH�={�(`�MD�<��D�!Dր�ja ]K����Zi�<��F��&��UȔm�yΤXr��˟ F{��I3���Is}D�za✾ ~XB�I�G`(�I��B%r��Z�,�bB䉵zc���,�4�KGiK��B�ɀt�Xd���1U�p�uAǶ�DB�)� ��[�H�/&�!�Y�w3���@"Oj<�w�E��4�r�؟*ͮ��"O�(�Ê4*$	�q�@�Z��aO�E���N�#U���H>9�   >    :IZ@-�nkZ��&C�'ll\�0Oz+��AI��e���X�'iD��  ���3]S#��S�&�5"�   �	  �  *  �!  �*   �pA���D���\�'ll\�0BLz+��A	��e�2b��+!��/f�<�'����L�J��Je$O�c=�p8�o�j�h���'^^� r/\�p����̰C2�cre�����'���Ss��/���O�(�P�Q�)��?A�����?�����'�����k��s$(i7��C�:�*�dy�'޶dU�2?n (�*@?K.`	��{�O 2������k�OL�0�'�P]E��##A�cT�I�X���`W(b��3�N=�)N�]��Y�QA&Q����̍�!��I[���Yg��:ɬ��',��x�az���]�c����ħ&���j�*̣#<!�d�'K@!��-ܑbkh P�(נ��O�Fzʟ�Z@NNi��H���W���+7+7�6��mh��ą%��4��G����n�
z�x`��#+1O�����ܸ��I[ƀ!!��}�~�!���$K!J���,���S�O�.M���.:KQ���<���雖2�t��Vc�/zĂ�Z��N&�!���.���ې�ԄLWI�%���#=�,�P-�?Y�Iʑ3|��C�I&'���.Lߟ��3h҂��'���y��4�БSG�K�1��夔?`A�L��];(���*=hY/=UeHٚ���yҤ̻r�<�(��JRWF�P �H��OR���?���hPiC�q�X�0R���WS!�$�<NܸAcS�b��q��L^h�⪴>��I���K>�l�L�/$m�l!�-��o �����|0���G�'�b�'\R��/\h@�
��'6�d>N�\����?Jtp0d�G�_��ySb�,H��-��,�N�(S֍t"�z�G��\e��C�"J�]ДD��{�U��&\]�Yҫ���8����/�q4�N�,&����O|l�ޟ̕'�r��]�84d�rƭ݁i��QJK�c�铇�OPL&�Ȓ�ϔ4�`c1���S ��0� ����%6�8��i��I5\�a���؟�n>^�0�9dʍ�f�X|b�+�w(�4��7��I�i��x�����`�Щ�Sč#����aX<��<A��Dg��O�<�Q�kE^�PڟHQ��`#�'֎�����?��O�Q�0�H�K�4�ӧ
�ZBa�d�O,���OD��?a���W`t-qbZ%DMx��"��	�HO�� K� �`��D�D��9���S�1��#� Ο��' �������Eڎ����ֈ�>Y����/�	�Tp�
^���ɞ$hpLY�ɕ��O]�'c"��2-H�|0Ŭ1z��ۅ$<�ēS��b?)DD�%\?r�ֈ�z1��ڲd4�đ+}�'��O��O���`2%#@�i��1���D<,O�9����)�cAN��:�v� �*��������'D���!�l/z���=xJ��"87iD��O��
6D�{���O���O����5K.�9e(��_��Y� �T7
A�^:>� ��6��D�Ԭ�fe�0v,%��?�L�8K������VM!�>}RA˓;����	}��E��	�6�������&���ݢ�r��`���p�2�(�l�x,
�i���'"!�U�����'��'�r�ic�Q��M�$G*ɚ���3|ܢ�I1�;�El�T�?y��7kh�!�4$�=-�\I+���ȟ��'a,�Y�'e�t��O����'	��"� �ȶ�ێ'ʞQqQ�ٖ)�@�7*{UN� �¯J즙H �>!�"�3#Z���Jˎ �6�JQ��2ʭ��� 5�1 "of�Ȗ#�:d$�Z<U΍ �dU�IJ�_�H"7�J4�:����p?���܊A��T@��b��D�[��@�L>�MSn��%�0©0$ĨX�e�Rܓm�v��J>�Q�[m�|�	�a+�%W��`�WЋ8#|�)�6�?������c�[�?Y��W� ���'�*���M{���vX�H5a��D���LX��u�����-K:-,iZ�2x��eKԹinH|:�˙���<$�B�`����M�޴l��Y�J�=�AS�*�]dVq�FZ�<��o��|rM<!&�W�u
$M�29E�����[�Z�6!p� *R2X��K�O�n�!e���?�.O�����Ŧ��矤�O%07�xӄ0·N�FqdL�f��-�lyZ�@\������A^��ڳ�:ZpH����`ӒO�,��P�F�Q�Oѹ]e8H ��R'pOl��#.�-yB���̚ O�;'mA�0��O�9�X�E��ݙ`C�&_�M<�#������I#�M#���S����ڇi��υ&v�$	�g#��qO��%,O�q� �BT�%��jHT�2hQ�:ғ���W�@�.7�'�Î;�p�бm��0	�M�R�W�Y�p����v�,���4���Mc���?������  ��'W�~E�ݢ i�#U�ѠgY<$��'����F&C'8F{���Tq����!F����IU�r�q��>aEo�>*���'�X�ɕ
av�˶�ZJT��!�O��d�O|�B�Oq���ߦY�!�;UF"T�;i:DQ�₅��xr
�G
6�8�C�sxmp�g��?� 5O��Z���ú���'���9S��P"���܅ʧ�UsF���
��s/0�)��?�����$5H����v>��!�L#jWP����Dl��hD�,Z �3g�)����4HfZ����>��5��eN�'bV��'Y2|��
��'�����w����OʮlX
L�re�*�?��i��7m�O�ʓ�?��}�Ǜ>J� T"Soԟ"�4��G����=	�|R��NB\�;�끗+��jce�Ը'�������yFa�;�?�ߴ:p\�҇��LlH;�	='0�0�c�'m�4r%@����'F�ɐ|��\PC���D �a������Y�.)
����٣�ay��H�b8qO�-�aO D6��p/��;�(�ش�'�n���wv�&Bs�6��;~h���>����G�O�x�'����	�Y"D���Sd�&	`M5 ��O\Gz��Z5	�0�Z}	��Bf��*�ގ�~�]�@!��:���������O\6MnӞ���V�k����-A{�ډB���㟤�ɵ�Ԥs���(��ҧbL<���L;f�n�"� ��t���h≞=c�#<�~�O�,�`[�l[:�ҙ�ÁJa�6t�����OL��O�c?����.Yk:��[i:�̲�j0�I񟰇��-�ȡJQ�Pc���&D*G�`|Gzb֟�)��$��A`5��O�;���!���vL�����O����O�3���ɦ�	����f}k�>~�K��*N��P�@��
���>�CG��`t�Y�!ړh��<"l�Q����a|a�-F��	;*O&(Ï�L<I�`�J_d�a0%`������tur�'!"j��Yh��,O6-�7,��Q��V2;���#��2`����h���Z稉1�|K�d��"F�	�y"cރ�O��ݭ�?��OĈVT�J����5u}��Aw�O`mڅ4���f�B�u�'� ������B��Y�`Bbxd�X�'�b���n�R�]�`)Z(I���X
�'�J!�!����Y�&�6=� ��qO�u�J�u���P�o�?�
�6�{�0��ݦ?v$�v�X�0EȔ�u��Oh�=!T*7�˝�$~pv�1��p�pAĉ��'����<�!�Y~��>�����_�f�b��@��C�	.;��@��T�:�Vm�R��CL�C�ɞB�j�r�I�P9�A/\�NB�;?���K��v���`�(b���?�Y2��?5��;���מ]��ĂE�'7���2��)7�)�&a�2uRG�̢K[�@���*"=c��)5m*X�q��'��1�DE�'��i��+_[�-
�'ڄ)ʥ'
2Yp���q X��Չ�yB�)�әS��aScY$L&�����gdB�ɍ5W̗����˗��� �:���&4���Ɂd�P�ő��o���0%�Тy��1�	%)�>�y2c�����!�F����>\��4���xͱ��'B�8Q�P�}@�����8ܦ 
�'�PHA�	=)?����D�:*�&iщ�$-<O1`FS�h���ʇN���C"O�(xB�!�����S:аf�'70�iё���<4K�:yue�S-��vḄH&��J?�7�i*������\��O߂0��:,ܢ��C`A�0{j��c�N� HdV^ �Ϳv+0D� V���q����კ$M�:gL�Ph<a�!G�d[
�H&D�W�C�F�[���#N>�EHH9O�6��ԋ�B��e�!�Z��hO��JLR���f\��8��	}r���d����'�T�<���`��S5��c3�e�A���S�Wc�B�	<i8r�2�Qe�]�$��?	ix��/��4g��-�%�[��X	X�\^�ZB�	�t(��ؗ}J�W&��DP⟨���?�bǙ�Y(�$���j�`$HW,�hOt�s�S̓J�t�� P|�ǂ���(�1I��	���@v̓}��P��<�3�� l�#�B���bҁ��=`Xhx�"O>���P>{�����B&hx�$��#�Ş<�&!Y���A�>0����D[<���OC�d�lɌ*�zx��
��z�Ќ��|����ے3�d��T#D���`��o�+v{RC�'2ʼc���S��O��M�� �84�'`��H6��� ������oX��a�	�&Fr8󇖂Nr!��,�<;%���(~U�E��
��؄牋+l����C�O�!r5$�2��B�I(l��!WH1Yg����?J�Z�ăx}��(���'��Q2{���]2r�+�@I?q��in&ب���O���7'I��9ڔ��s(�QH���[oh܂bO�=w3��
�k� _zU�� ʲ��S�X�|���P�E4t���
�'L`�`K_+T_
�D \�Y�`�x�l��'���k�IO&_�ޕs$H�9�V �r�i�Q�%�OVY�Ӏ��~����� �*���D	���'�\��O~r�\�� ������ځ�ϝ�yr�D�S� �Sv�X\�dp2����0=��O��pr�	�w,S&S,�0�lI>�y�o�z��.;�8�x�`��',x"=�O�V��@����S�G�39#�Y���ɮy���y����|R��<$�ɣ�bĜ>|8�§V���''�P��RR�g�1���W��5s�8Q���^��B�IK�4(�#�#-T�Ta���0U�:b�XE{���ɝ�O��]@�&G A^�����"�y2b��P l���=خ�j"G͞̑�d�O'.�p����MȂ���;�*���O�1s&+_S̓aG£|��EО1S�k�+<���`�['[��)Q���G����e.J'a�||�Q-�d�T����6D���5h�*[��q���R�T�X�"���<!Tb��	;<5a��Y'���p��}�<�g�zn"l��_;�*!�K����:�O<qDz��χ%�DP��a��,n,C6/QH���Qڦ��79�k�$�OTEӢ���}�-`�j۳"�	a"ON��#Or��Pbq`J��R� E"Oz(B��5(h�x�b���)�u�%4�Д�E+'��l3��6�R�!|O��&��s�0g}N`�.�#7�J��#";��]��u7��	�?���R�^*a史s�(���x�r�b����:��8�t��
<6��\�WѥG�!�$
�C)��)�&�3D�i��S�1�azb�d��d��&�!*<J�VK	�M!!�dI� q��A��7P�D|)�g=]��OUFzʟ�P�DkW ��I���%/��B	>ړ;��,!��¼��4��fJ�� �Jڤb�2(X�烫Pi1Or}�b��&����PU��1��&��HSQh�)k�Ј��M��T���O/g;F�����-WeV%�<����	˽k�t��`���,�C�K�v�!�$�w�X��Ƨą �j�1��Ϥ8�"=�,���?1�P�fo�xD��� ��q`��pk�T��'�>pG���������>������6I
]p�H�4��?ѣ��o�8�酸1nZ4X1��A�<I֥��P������S3%ˬ�C�
�c�'I�yR�
�t3�D��[����6��3�y��)��# �I=Q�:��臘�?Y�S�d��D�G��b���9uܨ2
8��� u�j����M�L_l�g°�{K>���'�~�Yf��'�
��_�<I��I�Zi�X'��41d��1���Y�<��� �Ԉ��4��玔��xY�o�r �1É~y�yq��M���=р�|��ǥ'2��)&�i�
ѺFCL���'ў���I��?0J�.v/�T���B�%.����	Q��b��84�,��
%x��� ��1�eN�(F�!�� �pA�@H/H����R�=��x��'��O����*�+��qH��L�N��xa"O�\��ðc} �wm�WF��!��$�{���)gN�bO�2OZt�.L�x�d�=�A%�?,C1O�"��O�DY��Um�Hj� ̯S�X	P��϶"[X�`��L>����/9���т�,WބɒS�<�灕
���pM'-��!�N�R��hO1�
��uG�	q�9��'݉7>�ir"O�4��wW�u�ר@(M1  �/:ғ��I�U�jF, #+��4B�8�ň�<z 5�	40Mܕ��y҇t�O^0X0��� Aڥ���JA:×�&P�t���Aۀ�A��P v�I��k��^��E��V->��@�Ǣsa�k���r뚄Ex�'������Źj��($-�W��i��'�b�@�%g�육��Y�UM�����g>�I��HO� &�@1��W&���I6��yP�	��ԓ�4r`���?9A�����e��!G�=� 1�@V/`R,%�ȓBz$ay � �9D�$�fB>�8�ȓE���8鍕33:��_ IH	�'aZqȂ���%p��U@9�"���q��'-�1�PJ��v�h��%H�|��j����
$%�ȓ�7��i�g煡\�l[D�VGH�>��`#�I�9�������Q*��cf���J�(R
�:q"O����ޛ!٠,��ŨX���ӷ�'��O�Y[���y�n�Cf^�J/���c"OP��7��n,0/V�{�6����d�Z���)B��Xѹ�%O'S-��PB��ZW|�=Q���)�1Ob��F�O����Q8^�ͳv��y��r��$D��PJ��L>!�"�O����A�*��:4pĆ����/Y����s�Z�I�Di�<ٌ��i�B���
3��\�8���'��?�!�H�}/t�./�hh�1�����	r�	&�	�6I.pAGd�F�@�ӊ�w�,��G���D�<a����pd�Fn#1�t|�3�6W���P3aV�u�6!�3�'�A����-}����[&���B�'Ղ<�EV;^�A v��P$��'�x��GL�7)p|i�H���'6���&@��L9���ovP�3��u���%�HO�$�8��H !�X�b�?
��V䵟��4*���<�g�*g�t$���$�ȬK �,ht%ǆ<�@��eL1D�ب�0*�`�QH	�"��8�m.D���+�n\�fL�
G��9dlC�	�;��8����r�&u�㛣kڨ��d�G�8Pe�p�K )J !2�C�+@��C��γ?�,u�I8s�b�p�hKR��H��
�\ft�'�j�����'��L~JRL�(&��Sp���6DJ\���s�<Y�G�[�Đ���m�;��T����?��Y),Z�D��M�-m�RY�<�4h�<ruHi����p���f�R��0Z���\�VC���Z40Xa` 	�CZ�Z��dV*j8�9�<�W��?Q��lό�lLȤ"�<�� v
L�W���"�E(�3�Ĝ<i���-_&~�|[��8!�d�d�����49��E�eʗj�1O~�=�|҅N���L� @ʤ+W�pCQ`�<��k�4��;�[ uZ>#�3�HO�ʧuD�Oء�s`�Bz̓�&�>�� ���'ex��sO8�	�MG��J,��	�ph��7���[�e1#�Y��E���?ф`X')���[2@18���@�^K�<���O0羌�g@�a������N�'��yO�.|m�D����	�<��y�m�)��I`mJ0%��M�6oC�?��U�h���D	r�ɉRb��J�(S�+���yB(Φa��	�C��Zb�1�I�C���o!�$W��$��vf��Q���S� "je!� [�� hf�NZ���`���.G!�� ��
4h�}� ��#`(|�f�)4�Y�j�$0�4L1��<Tyl�qQ
&|Ov($�����7[�.X�g�V'�⽈c�8�	H��u�(���?YL̃-�&	��]�����ƫ�j�0-�c����.��ط*�H�9dd�I��sP�¾?�!��Hz>$��ƍ%xr�u��M?�azb�dU%D���(wV8����Ų:�!� �hj����׻&��1�1��d`�O,�Fzʟ8�ӕ��o��ba��(Ve8�FL<ړ���zR�$��g�P妁qvD�w
�Uq��y"1O�W�E����MET�!d���!���[6,9�̆ȓ����0'B�d���XR28�<!���I�"̆I�r�<,��h��K�X�!�Dg�R��&MV�Y��1���.�#=�-�y�?Q�#uS��23,��[����Q�I>c8�����?A��6����iC2�'���'�NЫ��a��){��݉|8*�H���YnF�+b+�j}RK�J�dL
P�B��xdO�6�r�)�M2}D��S���&`(\i����Tdt���~&�Z���&U/X�j���2��$'��?��O*i������鉆>ѸhBM߿'m�<8%+�"qDC�I� �а�Do��Q��XcoKJ���$�<��L��
��'���T���d�9%7|�,D�d��͈�$ٛ��'��'��	�%"�����(���Y1�i�}1¸����Qab/��t��8sԥ�3.�FY��)g��1��
3�t<�`r:V	�֪.�b51��Ɉ(�5Q��'S���r%��QC�ȓ��BU��Y�<���hO�c�����Y3l;�  Lɱ ��t�=|O��'��b`,D?h<�E�`J"v��ˡ-!�ɴD���	WyOG�W��`�O_��N�)$`p���N��}���y#j{�D��O�ؘ.��H#6�Dh>���	�9~`xB�M�3a�X,>4�zckS�6`	T)�%W�xB�0y����#�4.�N�IĆ�\0���#K�4/6Wʮ6��l���'8����?y�O�<㡦36�*D�FR0|��1�D lO h�T�	4|�	r&�nd����g����Dq *��A*�) VT�B%Fd���O��j�x�1L�?m��A�$�Ԫ;��_�w6mV
SK ���RW��d�O��I��H�g�����3���O/d�B��K��T�ΥV0Ys��B#L78�jdM�a�q��#�*3Sרh����ƄC�,IIw�q�����<;��'�����?	���bӈ�[��U5. 8�H�5���"O���֌Tdަ0�4�!҈����$ғ������'�n�A��6A9�,� e�N���F�\�<t���OV��E1OՒ��u(�� �$�O~�	�^\���!���&��|/$	`��K�#�oU��e_A���Օ~&���gkJv��!�fcY$۶�Z�Ϗ�J��$H4�R�]Q��6A� b?O��� �X����d j�Y��@ԟl�'�6x���|R����d=d�R��tH@X:7A�#C�!�d �d�q��F��>��؊���f��e�4DM'��?]�����T�/����2�(Ŷ�#t�
6�JI� �$ya��������ПHZN:����	�|Z��P9{��I	1jH1sظQ���z��1�Dl\�#��B��'�V!c�ٶ䮝p2Z+:���=�$ ���{j^4�����3`#RL�
M 'sV=�@a�֟���M�'0�O��2Fccb�*5���t�'��O��#j�������'YX����$_,G�D�d>�Ir��Y��L�`��	��8�����j�ij��OR	��U/�1O|pʰ���`ަv)��/U�ZH2tL��y�@(�yA#�˚5*�x���ͻ�0=a��b� =��M�6���%>�xa���y"��;y<��FlJ� <p��0f���'�#=�O;z�(��U:Ef�|���I#u����=�IW�i
 󄖜Kv�(I�Y��H%�(J7�N�~�1O|�jd�N�ȸ��=sd5�@�E&VN=a��uF x��
"��Ś�Ĉ�`R���G���<a���IJ�r2�x{���1$���哰<M!�dY�fĈ��Đ�h�͈fd��G�""=i*����?�a+0Fju"b�Zq���hf'��<���p1�  @�?   |   Ĵ���	��Z(�GI�:G��8�d�@}"�ײK*<ac�ʄ��I&`�rLx��l�Ԙmڟ3�	��b�WÖ���G�,�4�شC���@u�I�>~��A��k���e&Wk�y��4�#<�o��q���*� �D�Ο`���_�[`C7Y}��#��$?'��nM 7-�i}b
3(h��p��9m�D��p��l����ƽG����J�<�5�.h��c��O8�,RS�I�"��1y3�48��5RdHHz�Q X,�R�t��i�	����<� %�Py�(��@F1|��U:�P�mv��'�r  q��'`�`�G���Y����O ��UMܾ�M�2��0�P�˃g��Q����J��!z��{���(x0�hUH]� i�)����>����_=�O��S������� �	h�Zc8e�h2S��h���"<��&�	'r� ��.Q��R�M�f7- �O6����d�k�X=��W�H�����׽{�XQ2����OP#�O�tʱ��5��5�Y�9t��Y�|Y&�	�/4�O�<(�[QRxx���T�
��D���O�܂��D��?A������5�HG9`0sAC̓89�"<9�8�	&g��HaFRWЅ07�60���X:�O��H<��]-05�&%=1<=h`�	��lLB�1R"9c��yVd�(�-�=vm��A�j��?���i&(�E�͏�?���";�����#G�`q�!kJWy2e�,��y⇎��\$��[�`� "c:0��iS����n�8"L��3�i?ʓ�"<	 ��5z�Y�ׁ�&u�(�9�@�<y��] 2  �����T����*v�!�DW;�F�� �B_�M�և�2���G���Z�0�+�BP�%Kn�! C��yrdJ%.� i��&>�(R� ��y"!�-}��I�m�	QGcī���y2�ɵ>Q �PP��},:5J�� !�yRn�y6��2g\���)#u,���y2��h�)��"	R�|*�!�yB�[�ZtL�$�v5��"(X�y��Y!n�{q����BU��y"�B"E��1�BCU�x�2E�0�HO
�񄌔�v�`ޫ\H
dꑂ�-n�����O����΃q��RA���h���u"OH8袤�#�K�9�F��D˻�y��.%��3��1 g��b嘘�y2�L�^���bCBZ*+V�a`1 Z��y��	   >    :IZ@-�nkZ��&C�'ll\�0Oz+��AI��e���X�'iD��  ���jZ(C�zd8�4o��I   x   Ĵ���	��Z8�Fi@�*x��8�d�@}"�ײK*<ac�ʄ��I&`�rLx��j�ЙmZ8d��"᭓ ���iU@ӂi���43�v�c��	� i�Y*���T:�@�cF�P�A�F#7�,#<I�&`Әmk��,ީswG�Z������$t�24cQ� $�	�N�z8ɳ�i��4�I��'�;4� ��V��@����b[�*~�Aӌ��s@b�ɵg�x�� ��7��8�
 ���'�u+R�/
Y��:��[%!����DP;Uè�*#k�{�剫f$$�r̝�P�)���~�YI>Yp��4Dk?�$, \L�s�m~����dlZ��$�=/����%���tġ�/O8��d��O�,ȏ�$�Gʹ�R-_
>?�t)Ţ>/1^!Dx*T�'B9�'i&�DO�ANZ���Uu�L�*O�H���I,i�qO2�[� �Pj�!j�7/���H�i���Gx2�l�'�&,�e��5qR��pM+I������'� 9Dx"��_~Ҋ+�lk�b�G/���R`����D�
�OHȡ�r,6�J��Z�=m��У�j8"�Fx��[�'�V�	��b�ͨ}1,iP�FQ,r�$���N��O.�qJ<�gd�
f�6�8
Ɩr�
<ٳ��k?��a9�Ob�zU@����P.K劽!��åPW ��Q�iE����Ο| �J�}�J7�H��?��iޘ9_����ϛ)~w���B��u\f`q��Elyr"[��y��.]�*�&�@gD�0��02���|����\�G 3ʓ�"<q�k�V�
�Bkƽ��13���]�<RcA 2  ��ʂ"O\�%�KfȌ�s$D?Zྨp�"O����N
%9:-$����"O� "!��ls���O�|��"O���*
��ڹ����>}�b�"O8Er�:��B
�x��,�"O��a��F�;h⑀g��#��T��"O>ȳ��
)��u�
޺D~�T�"O�	�U�L<:
 �㈇z}���"Od�W�h��)�(^�omZe@"O�z�� �%X��1/s�[�"Ob��wk�^��Q��S�U����P"O"�P��:1�Z �C�S�=}$ "O��c�d��H5�L�!�Nwt��p"O����d "T/ఐϜ�,�ʴ�"O60��獵*����$(�ȷ"O@�3B�@$g�͸0O��tyVe٤"O\�   >    :IZ@-�nkZ��&C�'ll\�0Oz+��AI��e���X�'iD��  ���4>J\�`"OP����   s   Ĵ���	��Z@��wc��:6�,0P�H��R�
O�ظ2a$��	���ī���M�Јhz��5g��@��9lK#��Fea�b�m!��=�&��jWJ�h����%�P;/���ExʖL�'B%mZ,\gf�(R�{�x8$��7j-�˓��C��rؘ��'44@��ަq3�O���� K�f8�(��V�~�R�\�z(fb��d}!�'.M�2@�<f�6���|B�M��DE3�KW�Ys�q�֏�".���(�"D4D�@˓v�4I����\��'E˞�;l���♡UQ����C�X����!Sh/0�q�'�8UY�a�#M��P;�O:D��W@`��0�'�@�����7�@0W�J�e]~�ɜ'�}Dx�^�'����ᗖJ]2i���!B�<�t�2�8��#<��>� �[��H+�́�I[�X
�L����O����{"���ES�-�$럾��	X�Ջ�M˱�59�"<�6�7L�Z��#j�+4Hٔ2�
��>�1E3�>5X�M�ͻ�A�A"<`k$GO*r���'�uGx"O_��P6p�Ң�6�U�$/ѣ7��P�b�(^�#<�"�Ob��c�~i��j7�(
T��Zv�$��O$�J<� i���R�[7:��(!h�E?��`(e6�O�d���1�١��hL��f&X�w���Q��i�1����� SN ��i�=�I��McV�3tw����
��t��& �<���+_M�<ʓ}�ص�1G�{�kz���Ո(�&`ʴ8�#�^�>� �	��!dG�G�Q��y�ቆ&���r�.���H��	�C�I%2�� �  �&��� ���{B��\�<� �1�te��RYj��h]�Y�(�� "O�x9S�2<�v�X��؜,���5"O�]� (ӑD���7L��w܈�"OR]�UHf��5yGՄr�r�I6"O^�����-���wl��K�V��"ODG�)�JE�%	[�6H�	�"O�P����8Z��'' +?�D`��"O�q�%��/���:T$�
~�lC�"OL5�(^�q��� W��Uؤ��"O��I��i�T�X&@Ȍ?�V��"Op��gLH:p��oY0;��q�"O�d�6�Q&jo����уu��"O�T���.!���+u�ڻx�!;"O̵��*��[a4�)���4�Z=B�"O���"��=^. d��%�v��Dx�"O�x�p"��*�8�$   >    :IZ@-�nkZ��&C�'ll\�0Oz+��AI��e���X�'iD��  ����O�M߸�z4D�2��   v   Ĵ���	��Z@�FI>M��8�d�@}"�ײK*<ac�ʄ��I&`�rLx��O�6�_.;��}�0��XT"![�e�w��n�M�Ʋi�����n�|��E�]3Q���ٖ+N+@�t��ɧn#���$�i����W/U�>[�M8�ŢVq�)O��ʑȃZݹ���I��Xכ6��>A�����x*U��:<�E��Ȕ�Z�4���R�B�3�{� ��9+��<u:O��M~�;��6?&��2��Vz.!��i
)ra�Q#+O��ĩ�l�Ƚ)�\������)h�Xs��� �V�{���0�R�X�&r�����l:H�I�j8�81�'9n8q�l���"�Ou+E*P��ÇkZ��h@;O�䙏�d��O�lYR�(G
�\s�a؞q4,�Q,X@�'̊�DxB��NyB�� Fbܜ)%j��g�T9p!�}��ˠ�O�t�{�Y"[7�$c�O��\�F�(�M�c9v�"<�7#Qu#V}�,�7FΖ� �͈C2�]�>��"/��� �VUb��R���8Q�擊n�:I�'�20Ex�Ɣy���`�F6��(��X�`C4��g /*��#<)W%�O0�h��>F�xтG.:؀�$�dX��O�3J<Q�^�V�J��#GDo�	�1��h?�P� �)�O��5��B[5 bƉ88 ����p��]�F�i�85�`m���x��'h/(6M'�?���i�n��Do����Zǎ�'��HXT�X�p7���$�EHy��YWv½��y"!MQ�>$'���n�(UN�ڧ�א ����Þo��	�*(ʓA�|#<aw�S�A{�� p�Ϊ8�i�C�G�<y���) 2  ������*�ax� ��Ji{&n�Z�nD�C�8s4�nT7e���5�F[4~�s_w�^�se��@�`]��v�<8 lE�g�\�s�ӳ�d=�m�"<��P��y8�����N�S�젦C�z�Z��Ǯ&���R��1���� .Q�h�
b.��+_��9n�!|~
�e+F�#���ҥ�<!�k�0g��e����>#)�]ibb�������oɘ�sFlҼmX|1�7ą�.FTԺ֌y�2�4#���G� Dg�l��M��8�V��O��z�FhFH4_�6���_��4J@�?��6�~J���.<� �d4]-jA��C�0��LaA"�QH�L�B�-5�-;A&2�8��˵^*fU����{�Nu>��ɧ�܌@մ�3HL
E��ɹ��A���   >    :IZ@-�nkZ��&C�'ll\�0Oz+��AI��e���X�'iD��  ���\s@� `�����oD�{�X��3t�d+ɞ�ui��"p�HRnax"f�K��{�NW�;G&���%�Pb�m`�BZ���=���ߜ,U"�Q�F�#!��@�ޠ)3����R�Wb�qX��(���(a��M���Ҝ��_&urY�?�D �	�Y��Dl�	Q䞽I��򠁟'j.m��ǖj�V��a�QT �P$V�bD���(<dM!��!}"M[J�'�uxD�نVbT�X" ޲.���@߇FV��ɍ$�9_�<�` ��DS�]���#�1��.���/ ��#U5A %�4��2+x(X��>A��f�%`��!����^Vl����z���]�R$k ,��(�Tȱ�/?n����D�Ê��}���YcEpM��N��;l�� �,RF ��hٽ鬑0�'��|�
υPl�iЋV	����3w��H`E��b��0�Y�>~8I�JTd�Q�k���䩟��S�"�\�1aH�Lf��k��,\ONB�C�.��l+ïT�LV���ƌ ,����f�ސ��2�]_d�҂�i�a|
� X" �O�t���Â�$�����2]1d8�t���9�Z�:ы\%J�	f>��k�;Y�K#�O#F`ؐ"D��P'���S������Q>�n��@�B�u��)%OZ�(g
�Я���]�ϿS&b�`�z�u@��Ȕ`���E�<1�eY�&��E� DTWȐ����t}R- ���"FD�+����O���с�6^fx��N$U���`�'�<f�F�p���B��)?��=����I�ؙZ��Jjy��'FX�I�W�|�5+U.��v�p�Ɍ��l�ɣը�,@�Nӧ�caE�u�BŪ�A�l�ಕ%X^�<!��� ��-R�'��;�0�c�X[?�f���8kp���0?	P�|�L|
��Z!J�j��5��B�I�����`h��fv�4�W�
�e��O� YrO�X��y��O��4�L=C��Z�byg��(Z����I�lԍRV��g�������6b���n��(i��/���퓮f��U:e�ӆA�h�{�n�;W�>�?�v��Nc?�a����m�k!Y�s2m��'��M���`,�R�b>�O.�է �꼳ċ~qv����>qw�7�S��u�4�PF�!i<Q�G��;ݠ����~Ri_y؞��g�ݙ �$��"S#q�r�:5m<�X��c���q��7��*���э}0�yz��U9\�Ɠ(�T��bń/��� �cZ��Jl��j5�	I?�b/%ҧM#�@���.~��4y���5�Ն�F����nM�MK��H$m�E�j��'L6)Ey����e�!'�0A�!t3�٢��$���(O1�p�R�%(i������1zV�=��"On�kF���E���(¤6����"OV��ÊSsଁ�&O-��YPB
OD�iŋ�'x���	��?����Y �y��_�@�m�3��aQ�I����<Q�;�	.h7��J��
^urɓ�X�?C�I��܌ɵÀ-�X���oY1s�>�OZ�ʎ��i �ɛ�k�,��<�Qk$,!�$�-]����ꇞ~`֬Q�M=��!��'����^�z�8���G�%JX ��	�'sT�䒹Y4�bn�"KL�Q2g �L@,��U�
!��-�Ԥ�Y8�xm�'�2L��D�M���P!+D�|��
0l7���!�$�2n�7`���D+,#P	��A�>�J�E "��z�b,O�P}��Ǵ�?��c#zP�	��Z.n
J��e�i�<��c�G���"ˈ."szd��)BN�'_~�GGˬ#����F]{���;V��h�*�&u�B�Ӷ"O��j#��2�``�	�2|d���"Of�cԂC�m��|C���	m��b�"OV�y���/9y�i2"�G�~I�
Oʴ�`�G!h,�ρ��ph�W�ۛH4a4�&�O�8ːH�"a�� ��M�2ʖyZ��'����=i���O"��R ��,��6`���J��Ol	�͘6�0>�	�("}��r��8�̱���EEy��M15Q�D���1��P���>��� ����-G�X���b�K!�(_Rt�"`�a^�qC��� f�0��U�p�� ����t
ו�� ßw�� �wJ؍h����CB�P��]h��G��(�'�YG~�yAf�h1��aȤoy桫uD��`��'�����	?-��~BJ	�&(����U�^�Du�F���O��H2�NR�P�C42Q��$	�XQ�э�q��� Ň�֟D���&�l�2W�'M�=�P��8(�tY7L��gAd(K+O�����33>�-��l-�)��68�9����M�w��3�(�,�1 ���O�x�<Q�B��U&�h�p�.�HE
�5!*��'Yʡ��T*Pь��V̕D�D�(W���]��3A�:�H��iƹI����$܅�pJ���	}���.ײ�Z�J�)�'��p\��ɎM.�g�y�̢Fc��K2jy҇�Ҷ���$O�T�kӿ����O����3V?��u�ܖa��`Ѕ�Ob9K��Q:^Q�e�ucV`�E�4xC�m��H ƕ�O4��[�B�O���ۓ�J�;��'��kVO·w��u�PE�\�y��'��t"��F;��` �H}�����<p��|*��� ���U���.%�M���%���4"OĉHJr�h��	�i��+P"O�J�ȇT��8$ #j253�"O�8���+.\��F$a>M[�"O���b��m�1Y��C���C�"O���&n��&��H+���#Y���Ѳ"O�se�܈�u:���̼q��"O\�*gK.�DB�!�:��p"O hR��A��4�����04"O���#-p��:d%(r��p�"O��(e�,/�,���M�l�Rw"OR���9�AY� ʺb�L�r"OfE �J	�Iy�)�^�"h�[2"O�%�qI��d�<pYU$QH�h�'"Oȍ�� ��x���*���=J�k�"O��A$��(?̄1���n�	��*OP����z*z�K�D# $�S�'��Q1�Js�ҀR���tF�1q	�'��p�k�&,A�%X�hU(�A	�'M\�#�AO���1S��euF8��'lR�pG.$Y�e)�n!7j�(�''���@����eK�u��9�
�'yl)��©]��e��H�ve����'vĘ��*�,�J<�c��^���2�'fP��u�mW4:���D64$�'Za�ƈJ���Q1�6dY�q��'�"�@ ��8�*�EHMI�i�
�'�����B�/3�.6�J-c��YK�"O�q�.R/;��tbH��|ۆ"O�	4 _��|�� Q�>�ԡ��"Op�GG�@}�e W��&J�i�d"O�\K��6�.�r��ȋK�>U+�"O� ��D�Q�jp R�*q�b��"Ox0a�	 z���g���^�
�"O@�	w*+�Xxc�@�9�\#�'
�� ���7>��:�Jm���@te16É�h,Z���	��ȓe2��.��LoеxR�]*L$)�ȓm Ő��F���Q����V����ȓ�<PK�G3S��9�F��-�� �ȓS��mU?8��Lڒ�/z�t������=;R�0U(��z{���ȓN{r��=klz�!@l#be�ȓ^^4�E8m��4��^�����+P�Uӕ/�H�U!� ܨy�.H��v`h@ѩ_��)��I�*�`̅ȓqN��\Bz:�PAF9,W���7����N�"��� Qϟ;4�4���5���8��5wxEx��6V�1�ȓz���am�bZ̡��6]Z9��*��<yΚ�b��%@"�W�W��i��s���
��'�z@��
 �%
fp��p{X�I�HU��P$�T��e8D���(��{�V@���-q�� ��6D��PW�p.,���)C��!QK2D��#�W]�Rc���0~��ĥ1D�hza��K�\��%)ӏ���vk!�ް=U&��狛;�=���=^�!��N-A�^`0 Jr�,���m�!�
\�4�)�
ؖ?�y	�'�y!��\ _"� �d�e��m�EJ�9�!�D_�uB\@�蘫
%�p��
0!�ǍH�>��rjл?�l1�� c�!�[170�g@϶d�fq�e��9!!�� ��I�L�/�F��en	�;ﴍ)"O�5v�җcC�봠�]�ؙ�"OJ�Taݰ�t�"���E���3�"OJ��.�1l`��d� �����"O�� �g�<bfB��#l�E���Id"O�`1� Ů9:�)'�WO�H�8T"OHqP��R�t��E@��9W�*�{*OP��S��1$k��*B�Z
T��Y��'��4I�k�?r�0RB�G�#He��'-�VE�)�ޠP"Sg��=��'�L]!��cy��$�R�T���'�X��f��r��p`�D[;K�b�'��H��mC#����@<*����'�0���I\.Hj�h��fL4�
�'3ԅh�J�;6�m G�d���'J����M�P+�C�-S�$tJ�')	��Y���ص�ǾP+`���'��pQE$G:I�m[5��iJ�'�.���dS�t��@��W(T�<�`	�'�L���ǆ�L  Zj�a	�'Ķ#���>���r.I=!���h
�'��d�� H��q�JN2Si�P�	�'��<j���(j�����4�4���'��8$IA"T�=��j¯	����'_i��n̈;
"	���L,p��'Z��c&��v��� ]b�%H�G�h�<1��j Ũ��F' $rٛ���}�<�`��n��l�S#�'K�x�C�YP�<֣�\��A��;x�ċ�eM�<��DдG>
�X:��5dII�<���2o�ģ���2Oe~����TF�<�a�Z��vE."�.�����C�<Q�ز�f8{� :?XP)Í�|�<�.<W��U0EF~��b�	@�<a�L�ı7!L�r�Z��@�<a��F�8-`$m��o����V�<��#J( 2�:QNM�x<8$A'�Gy�<IrA���<p�m �o��ȒFy�<q���0��8ւ��)������w�<�0+��(*�2��I�<D�$B�#�z�<�Q.T��A�Ƒ+.]��Q����P�?�)��<�D �'h�T�r�B�S��K��NC�<�3�����*CJ��iȕ/��l�яJ+0�@��	���S�A* � �f��B\T��$×b��a"(��?Q��Y�H3C&�8l:�	f�E�<�T�ܸ|
1���@���	�{�|`�e�g�S�p���}rpş��H	�'�y�mADI�<yD5�B�UHG��)��ND�98#����I�H��	>P]R�q�W;?qP0ڶI�:���h� ��l�ax2�M�{�x�⇊U��\�O̱�M[%/��T�H�r�!8<OĴyu�7d��C����R/���Z!K�Rec`F;ON�`t�S1n�"�Z�#�`ct�S ($VD0!	�0ŀa#�Jv�d�$Yc�	���l��e2peD
$$�'��qB1���p�����Y�Z������V�l�yBg酙��O�<�0��ò#�D�Å�O,�&�r�bA��2<��>\�� *C/.�'�2�?�!�M,{�h��l6d'�m�T��������,��V�?��5�٬|R�Q��,Ŀl����0zc�if��9+h�cb�`!��O���A�ŗ!�V'?�XÔӊ]�9�*��$�J1ЗFsӶqj1+�2@;^�P6D�+��p���O��q�p��iڧh���)T�Z6�h`��2��u&�K�G2�m��� $����l�18_2.�6\0�3c�6ɞ��U��,�
D�@���a���ld`U��. ��Q�F�d��\n� ��D1z9�ҁy��1�"O�2c�HQ��� !P���	^`z���b�s�̹���{�2����>#"�iW����.z��6�� X#(qd-�Yi� ��V�T MF�4�(*��S����C2�x�����~� �3^�E*�b^�!���$�ʌg��<�O\q����qO�%���Nw�\ҀA��w���H�W���I�|���#��>!xw�<� �0�T#�G���`���.�K�AI�K7����ޜ5��5	I�>m� �]����i.�k?A�ɋ������O�@E'Rj̓jL���GK7I�)H��i����I?ђ��+
>pA{R�� )�ĤH���<^ڠ����&��}�m�2����\� H�P�V�T��ODdh@�Z:R)Ľ���%��� �ܹB#ĩe�@u��ű-g!���Y�g�8z���M+����3>����Q����)ڧf6(h���(f�@i�TC�O����2��V� 6"߮�L����O{�$?^c���0<1'�ČL���t����!�t�_I��T�'��?.� �#���u�*�$9ѢË =!��Z��Z��&`$Hm�ԏ]�Q���j�SDdp*f��?vt���Ç���D43�!��7F���sW�+k-�@��-[>4��d��y�Hq;!�¥��)�'>�ԛ"ͨ�������/�t8��J����A9f
���
�m��O0��W�U�j��,�JLʒ:�v��4`�Q������<"@M�U&�%6J���k�-E3R�@���da6,�]V�A Ξ		7r��P�E���FRD�8z$ ��~�RkA�n\�љ���]aL^�<q׃ǒ	|���E���+�[�<9�j,RO802���N�ތ`��XS�<���s*�\h#��&k�|�r$a�S�<q6M�0�$�ɏ&VH�3ft�<)�G_b� -3"Ŝ!u���CV|�<y��	4U�ƥiVf�3@$L %l�<ikl�9�C).y �:��n�<!�BO�P	��ֱ%w���$M�<���r&6�aD"�WP���M�<q��^)�*��'/٣B.�z���H�<i�(�`�y9�o�58T��OK�<�6�@4C� ʦoQ�%�l�j#	�M�<a%kڠw�t����b
جZ3��F�<�Q.L�k�F��C�"C+~�t��I�<!����A�[�AEA�<y��I�O��!赂ރa[� ���[B�<!`b����4�D6O���Nx�<q��ST�#k�?C�rJ��a�<�l��g���0C�@�����b�<��Eӻiˢ�Q�ʋ.s�F��E\�<Q��*��凁wY.���s�<ѵE!|�\�Ip��j*&-Sm�<ᕍշ,*�r���Dd���"j�<ɑX�f���g�6aI���j�N�<��m��C�N�K�@@-NԶQCC�Q�<1B�ܟFf���²B�Jl;$Vz�<A��hA(D�����TP��q�<��M�1�t�!	чF�	�Ds(<Ɇ��Y�n}��bDUb�+"&��GsL����V'��?A�G/I!�`��5a8LM��*b�xY����y{��q�>a���;4/ި���T�~�$Daei�b?q�.������&j< q؍,̒��%��"��	a2�,sFgW=0f��|B׽1f�����x�+�����|��*:'�z��ȓ!1�l*�_6���S঒�C�XZr�Hfyb��N�]г���#���O�5���s�9�­8�^�8�Ŏ*q��uI�'1�O-�b-�Z)2�
��  c��a�B�YȖY����*6D`J�$���D�Pf�$?�	4y����7KU�ȁj樀y[l�?��_.S:@�C�J٢��)N�r��,��  &���%$�>��j3\s0�\؞�@�hH)cZ
,���-�����䀣y�R��o��X�쓟N�Z�o�]��Pݴ=��Q�a�
*kB̻RcO��ZE��x2���M26E#��YJ�JP�GcYly2��b=6u+!���b��L�O~x���{ޭ�(�H�V�h���dR,H@��9�O��;�Ȇ�E��1�P��D��CpnER���	�U{I�Ԫ���&&?���f��B�
��9	���k�x�����V}n�a d���)� �]7��=A���ǃ[�BY<QQ6�'r��#�/�9�!�� rZ� ���J�r,�F��j�'�f�H�͎�49ɧR�N7=�(��V�$�r���r���w>@�P�"O�m)���I,���+Ό�f�b���-w;�W�n�OR�����[�vE��%K�7�8t��';�)�!��LY�$�q��';���U�R� ��
=�h��'r��:1�ֳA�UpRe�-z�|Y;�'�	j�T���E�Κ8f�!�'&��s�!ʡ��l����0P�0��'��EB`+�I�0B�U�%N���'4jm �GI(~$ �� ��*�'1��	B�� /�`�Єa>�x�z�'ց�V/�Sa��Tb�.}#*DI�'�DL�g_&A�!� Bh�2���'���(+(6u��u��54�����'�Ղ�d�Jހ���)6Έ�{�']��#K64��L��
	�"۲��'z�����;��5����/̑��'�pj�^��)���gq� �'��D�G�5O��"f싘X��q
�'�&���%׷0�R�e��9l�x��'��=B7�S#{��يj��l���'�T�Y�N�PLޙ�w��2���'�|@X`�3�,y��BX0\n��Y�'�6���^�pX�`E%�J3����'�ܹ��m]�t�*�@��::�x�;�'�4zs�lcH���'\�F�Ҵk�'g��� `�'z*0�#G@|t��'PJ�����M ��Z�2��|��'{$#7��R�(�Y�.��-~D���'����%��07ц��T)���@��'�FQS(�&�\�$��^~̹�'�v���S��D�c�C\�
:�p�'��ςil*K&
��N�z�'��!��3C�lY�E�J�^���P�'�zݰv(��������ʌK6"��	�'n4�c�23�ʥb��F	֡q	�'ˎ0v@J�{���c�%"���!	�'~� Zы��@��P6I�6��H	�'^Vas�K��0徬��%Z������'�������XUGE�f!v}��'�е�G.Q"�X�
0%�`���'S�E�E�y�����j�"1��7_N���-w>\q���=��q�--��0���`�1À�4�l�y�/���@T������vd�$�_��؄�EA4��
�|4 =a3&�8��`��Y��P���nq2��I�Z]�ȓ����X�'x��2O�~e�l�ȓ���C-T�Mt вE��lͅ�I���>"��92)�~����3�	� i���՛�G^� �d�G"F$����)J�5Ө�0�mY�@�X<��O�nf�PP#��<i�D<?к�E��ݟܩ���%��!�kt��(��<���_.u!ұ#�l
\>5q#�9%]�� V�Xҙ� mg��[�e�!`�C��)���S<B�h��3Ŏq�pc��rC�L� \0�e�bƺ�S>� ��ǝn�S�h�d��D���ŉpz��	Lyy�B��0|�B��4A����Mub���ꀃ.�xuAD��h���-V����8(���u�&���LÝV#���2OB�`B���~�6�a%�O_�u��!_@>�!a��s�I[��'�1	�#�&Xbt0w �4_�q���Č��(,�3E#>&1G̿�!�.#J����53e��
N!���,PqRL��a}����Q����"O�Xhl�9��ݒU$^/kp�20"O� �4�E�Ƶꊄ�t��^ j]�#"O��0���n(���ǙB���"OA��37���������.��"O097��w�\m{�+����*P"O��6���hJdj&I�8�D�c"O�e���)P�n8"��M�o�iR"O���7��T�����K�.��4S"OT�H'20��|�kL%O��Ԙ3"O��Q�B�f�6�����3����F"O��R�:}%���:��i�`"O�t���|Q��΅�7\�1��"O�,�Ҡ��Ag��T�]�9Dq�"OvIȓ��99
=(��8A��;�"OJm�$�I�����h��Z����"O\��D׹�.���MJ����"O����FpZ3���Tܴ키"OXh�$Ή�-�8+T�<����"O6�;g�$�,q���g�����"OҰQs+�14꠻w��D:rP�"OR�0s�*֭��ܠc'��cU"Ob���֦���HtH7	�`Hz5"O���f���J��Z���Cc"OVaRqI�K��@��͓N�H�c�"OV��`h\9�������-���B�"O"(����?�¬E�v9D"O`�Q獎u-�����|a��V"OL�y�/��%����I/[*}H"O�I;��ȸ&`��U!�206�+�"O�eK�MnT�� �дM\���"O�L�h�i�L 1۲s�@���"OxD[�ˉ/�P�+�F��	� ̛�"O��%��QQ��
��ϷM_v�(r"O��	9W�>��ʖ�',�
�"O�ђ�I43�fL�Vk��Q����"O�����M�s�0�3�l��|� �"O8{&a�!#!��ѕ�_/k����"Od���W�q���g� �	�hY�!"O�laTIPDjv�(5�L�;����"OZP3�h F܃v� ��"O���a̍C��h%R8J���x!"O�M�rg�K����rM�2����"O�Ѓ emO����/�Na�d"O��n	*T>|�qԾ\%�R"Oz{e��*~}��q��*� �"O`�0W��Fp�KE �8� ܹD"O�(���3[�m��nF
Q����"O����.�UKvt�ČX
iL�a�"O ���ˈ9
�gL��{���+�"O��b�e�<`�zVL��|�̈�"O�8Q��S��̐e�:w�e��"Ot@�FAD���x���n� �j"O��.������H�p���If"O�4#�C'�kZ)T�fU��"O-
�*T

�J0h�j�$6�U8�"O��f���(zԌC�V�?)R���"O���煗R4x���M�OВ�"O.a��d�=^��!��P�
]�E 4"O�E9ulQ�z׀��l�r�VH��"O&�&��|��i��j»e�Փ�"O�Ex�@�@��J�.en�e��"O8�����b��Z�	K6Q2 �c"O�mb��ă������#PR�s2"O��b .L&�8��4�Q3( "O4LS��9�Nl����_ �y�U"O� ���s�	o��Q�7�S�EPA�b"OZ��@�
��� �oE�`�Ve!u"O�<k�'؂��*Ġ�7�c"Ot��$̟�-�|M���؏�dd�"OJp�QN!jB��0�VU{�"O���cg��Nex�˟�7�ڗ"O�ܸ�P&3�8��	�g#�\�2"Orݘ��;	X�S"���q9��H4"O�=��f�2+�B�aCfL!QX�2�"OɊ��e6��r�nI:��\ic"O��@�Ʒ 8.����$�|�W"O�Lc�6$<�\	W�������"O���kFrϔt�D�f��Ⱥ"O�|�Ā�z
B@��+}ў���"O� W�G*��C� �:0в��"O0�閆������/���ԡ"OFE��T�qh"�T��!V/�4��"OZl��+�?@���Ư�8,q.\� "O��2��ʡ��w��,K1�`�b"O�)�*|�j��C��H��"O���eH��R�M'l���R"O$`�sM�:m+���B���S�"�{e"O�y�_�5�����%}\���"O ��!	�$�u�-R�u�x�`"O&�(E%�	5�j|���R�FưXD"Of4[�����+S�s��=b�"Oք:wO��>��M�P"h�*���"O�q�*Ū'���hfÝ6NK���@"OI;p� �s����Z<D�JT"O A��:|�Ґ `&�y��X��"OV�HR�y���! K=p&\��A"O~,"�o�{�����nQ+0&���'"O8���ΈP��`��7�,=�"O���P)ȱ$,����y����"O�ȐI\>0��!GL<�t�(E"O��p B�ͦ��5f^�;���2P"O u1��^UF� #EFȽp�R(��'��M+��D'Dޕ��oF�s�<���'E(P0Ch�5�|a��d�S�'Ap8b�/R,?�n��0��*[����'�MG�T6~1��i��D��9�'�*0c�Q4\	��B�kG�oKd0��'_���bX�oup;u&ޞj�B0
�'_DM����5dn�]��'M2�.�
�'��< ՙLP�dn�-y4M2	�'O>�����se�R�N�le�a��'�ӆ�Z ��9"N�b�I)�'�,�	���=I�L�j��BrLu��'n��!EO�m�X���R7G�2�'2���u�ˌ�~��l�7m!��
�'E�=��&� '@�QV��
�'�`�VU�{����,�;�� �	�')|Q�U�ԩ����S"#9�1�	�'�4ZWc�4j��Bv�I�D�
�'H��j񠚶y�0��l�':�<k
�'�x����%:~��hȳ10B�A
�'�x]B��	~¸��a�,a?V�3�'��l���H;Jad�[�%��YG�\��'���J���ij��G�cjj ��'{�k��Xh]�d*��b�<�s�'H0\��'��!n^<2Ċ�4#� (�'�\��A��=QP"4)4�ڨ'͘��'�:,�A��-��σ�#���i�'�t�q��S��C3f�7��:��� ����'#[8��J0t�j��F"O8�ҪA���y7H��^�BE��"O,%q���H�+(��!#"Ob`��-W5`�ȀU�7���G"O�����q�Т���LTI�"O�!�V��<���Tb�:&�6-�"O�x���$�S�@�&Iq��U"Otu!��*�	�R`��#�"OxyV�L�"�[3�R�xs����"O�e�K=�Ʃ؁�[�"��c�"O��6�T|�>��al�H�(	��"O$9�a�"��=;�*Q�b�n��"O�`6`^ Ͷ,; ��>xz m
5"O� �da�-o�4��i�*FD)�"O֤�B�Ң;h�m�N �Z.�(# "O�Eӕ�;X���է�73����"OqB����Jb�W�}�~��2"O2ͩ@ �B��D�ńX5c�`��!"O
�+'&�.g7��t#�7I����6"OD��D�n=y�����Õ"O���!+�ڰ�a�	(,�6E�!"On�B�g�(,Q��+��V�}1̀0�"O��Q2V�vᬨа,�A)��q�"ON��2A�!n8Yh�l�1kT �w"O��A#Ƈ(��Bá�)IN�P	"O ���Y6S��-W	�j�"OnQg�Q*_��;U�}�U�A�<��
�P΄�a,Rn�Z��0��~�<Y�^
a.�؂�]��E#��@~�<�Q $<���ZV������%bTa�<I��4`�Xd�E�?v��:TLO[�<�A�c��{$)���JtB�a�r�<��k��Sre[�c���zC�	��fq���a�T�K���
LVC�ga,� S�A��("�u�NC䉱
ߔH	 KՉ}V,Y�ҭU2$:C䉄I=b��ǒ^aQ&	R�/��C�ɄdX��
��ΫV>�EHC�l��C�ɋt�>UXӫ�z�0 ���Av�xC�7oH�C�J��ǌ1m�|C�ɋn��x��ډi�&�8A&�;=�B�I�P�
�X�̜<8���##L]�r�B�	.(���ȳc��	[~�T���2`�C�I0CV���)����`A���C��,V��u/�^����k<d�nC�I 7䔈(#�G/i�>ҠC��@C�ɯ\��Ui6j�?_�,\:rh�d.RB�I�W� xH3i�	��ūd����B䉲mB�q�v�ޛe����¬ �+}xB�l��u*� 0~���B��[E�FB�0Æm�'�3yb�0!�8	GC�I+`�vA�����a�b�;Di�B��X4���\�=P�����
H�B��>n�0\q`�E,&� �:G �a��C�I�Z!�ً���;B�*�R����C��=}��Cō��,�^�P"�!s¸C�m�<��$݀/�N(�+:��C�	�VarD��jC#D�GA �JC�
2�̔ؕ!�|�`�a �A��<C�	2^�\�b'���x�E̜�K��B�Ɂ{ ~��Q�}U*u�4
ُ:��B�	6e��� �0)�σ�Bo\C�I>.�~�� dӨ�:�j�,!nC�I�\_�P�@>��$z�F_A!RC�)� ��	��P�zQh!g\�XX:�" "O��؂̃@�Q���=a�Tt"O�]i�� ��)���2���1"O�{�G%?^j�
P� �J�{"O*� F�)Y�j��JcsL��"O��àe֒p�����¥oeQ�&"O�#Pn��dgt�Q��^T�uQ�'�nb�@�D5����`�^XE`
�'ҵqqm#U~|����8I�'�,H�   ��    b  1  r  �  "  D(  �)   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�H�!xn���G*W�(:h�.|&�t�BfE�C�V����5��8b��M�5P>D���@$K���x���1Hm�� ֡mD8�3�̕�Il2�"�JMz�8-�t99��'d5���!"ӫylhQsϒ�UT��VJ7Q&��&݅tΨA#�7z]Ҝ˴�USX�\8��!s��L�;u^"�z��9D�D�ҡ��[�z�{U���Й���*D�|!�*eZ�h7��K򺭁�*D�H�� z�.�ك/%��qu�:D���߅Mu� zBb�,5�f����5D��ڵ���?�i�d�R?R~�覬8D���RF�  hyI&h��D����&8D�P�gmܩS�d��wቀ`v!0w&8D�ܐu�lR���W+6�p��Sj2D������~(I���;�`5�#1D�h�ŇOB�t����Q�y>!05f=D��+!b;��)��p�X�(6�;D�8kC�|���^�gHP��6�<D��ʳn��v�Ȕ�-�IP=� <D��
�����P$�9v��!���y�B�9�~���,�zi�I �nފ�y����w^iZ�n[w 9f@H��y��Z3;+$L�RmT�7���h� 8�y¨�IFܳ��V8��&�ɹ�y"d�>xRLɋ�ˑ�Wj�ƌ���yi�$�����N��\�b������yr$�twj��0*e��Ā*	�'lp����=A��������=����'[ZԒ����􅛱��&;h��'-�@��Ш�D��)F�H9����'�@}���0c8L�F�
�A���	�'u��@K:ɀ��AF K�x��'by �,S��>$q�FX:�&x+�'�:�"��Rx�S��R.,�~���'�l��e�S�=���+��ܒ�'~v��锆P`�+��[ze��ɲ����w�^!A�!��lU�<��5��@x%�DY�T�ă>xa{RD"8 �����6+Tm���ӈO
hC��7!�b����p;a��u,��HaZ� �3�"\I�õ�ybBL:ւ�;i�<>*�Caÿ�yb)��s����᧚T��:bFD�MG��� c@� ���.����B"�
�y�$�^qp��N98�L({p(�=R��Y���M+�EO�E�E�?5��}�	4I�,X�k�U���5���0?A�, I�%�+x�|d-YC�����,Z���I�7p�Г7�'00Kg��>|+@�g�իE\کC���F���Ӆk4���{��C+U�^w��!œ[Qb� gb
2R4�2
�'�XXU�Úr�2D)���_N|��'E��(�-K�B^q���Ϫ��X �t�OH����Ip\�p	�m�)
�'�^���m��1���FL��D:�M�G�)+�F8ٴv�)9�L�i���7��'�d�j�"<���p5�ذdjΑ����I;'�]-���D@��Kl�C�!Bk�e`�旫nD�����F*D[a{R���ԥ����RN �k�ռ��O�}������PU��Qmb��U��uJ7HUC!MĴ[�!��L���y"Ƀ�#f:�I��=���R��o?1�ED�/lA�7耆j�����E���#}���ə��PA��|�n���U�<�A_8D!{�n�_�P��A.�&NPt��QE���PxHE�Ο��>��	�<g�0K��~���Ug���s��m�fʱ�(+�eiU␬8�r�`а<�Ή��fS�ve�ɻ�t ��I��V�0�$ҙC�D�F|���.��8�SӚ;�D;ql�8�M����P�e�����@/C4��Ņ��0e�$�E�r��D�[�7^���j�ܔ(�Jðm�>�y�@	+�eo:�'M �aQ6�J�[���c���.D2}��l��UЇ�͠_�f[2���z��	��LP]�ZoڼB�x�WK&���i�{d��#�%��Zs���|Q�0��I�:�"�5� ,��*Y	�z�Q���?x&Dz��� ~���2��	E����I�R��i����!
,ƉQ��/�4#>iSnW&mS|:F��(*�4��!������fhǯ"E��U��dM#�"C�ɟ'9^)��'�!�ؙ��X^牒x=��p��)a��Q��؏y�7�Ӽ:�@Cn[�����&�(��B�Ɂ�Fd��B�{w��z��˅���oL�o7�F��Pq�'R�d�6���5v�ѣ��ϿaT*�j�����@����|�D���P���<�T���Z� Q�B����xr�ēh\ yc�_؞p�'!�2�+�/P?`
���7����`Q��A�x�HI�C�|�oz�ey�2:%B(��(���(�l D�zP`F~���� <��H��n+D�� P8l�$�0�΂�s��`3Ŏ7D�XEӮ3X�	��d%��L��*6D�
�^�S�b�r�E��`�)�t�5D���jW1%�0	W$L�>��Emo/D�PQ�
5F}�; �����`/D�Xx�<���BfP���#+D��z��D�4>�B3�G�,��6D� �*�,08R9y5D 1{&H�@!D�����8T�z��lܥM$�y��.D��#��R#�̛����w��c�'D�T��:XQ���5}�*���:D��I�LǓB0j<�sU*���R��9D�x���U�<\Pvϖ�0b��J�M3D�(r拖=FLAI�*7*�x	I�2D�@�5��2Q0)�;ydc��>D�A�t�܀ƌ��o�ɉ�:D�Ԉd@�i�.83
[�Ӟ08��2D�$KO�(()�eڵ*�i.~�!�$х<��)��.�<9�d�f(�,u�!�$O�6��2%"��r�:8���;B1!�d�&j�2N##��\�-��!�ޅ9������;��V�D�F!�DQ0���C�q�j�4lϤ]!��5Ys�*)�P�e�N�
!�$�u��92���8H�E��'���!��s�r8���	�c(�je�6�!�D\<�R���4���p`���!���\��,Y�&	�b}��%GC?�!��C�z�}Cc�(ij\���ρQ�!���O�ܫ1��T���ۢ��."�!��K��"�Z&ʠ�nQx��ç�!��H�ΝRs�>X��Yc4�T'9o!�Ԥ�Ԣ�@G6a�(�<W�!�d�wX�Ce)tI�4�3�S!B�!�D�$6�%����m����l�!�D�"X��(R0�M;w{� (��<$�!�N<A���*R%D�&d�H�m��6�!���9t�F���d[�����!G�"�!�d��2���IJ�n=�Ac�g�2rv!�$ѠC�1`K7x(�ҳD�!�DV�8~��o��$�v�e�1L�!򤒱4k8�N�8渵�f�ƗN,!�D(�h��qʀ�*�RU8�� p!��B�|h:�A��@�<��`��!�D�q�v�(�M�M\v�'��!6�!�$��[P�t���t� ����4q�!��!&���FY>+����ç��i�!�d�5���0��b\�8��E�k�!��2 �󈘇7��%�r&��e�!�D�a��A�DUl�r����*(!���$�p� [�NcF͹r��@&!�d�*�J�u�$Xj��)*}!�$��@��s!��`���p!�� �y�`N��u�t�v@�!�H�"O8 �ΨN�L"�$�X�J�2�"O�a�o�"rӘ��A�	��3�"O�z���#8f�9Q莪(�JM�S"Oh����ɉY�v� .Y��F��"OF��u��; H|�pJ�਼I�"O�T��� n���zr�Z7]wn��"O�p��9{��m� l�r*��"OJ$���L�X�(m����A	�]��"O�l��J'Uqv�Q$��+���P"O�)�ʑ>
M&��
��h(<�b"O���kܙ.�FX�G
J1kjl�"O(�3��- C��uI�� P��r�"O��1� Q�Q����%��XK��H"OƠ�wF UW �@���)B��"Oj��Qlf��� ײR��+"O H[�B�8��@a�H@�e��9`"O^� �/�y���L�
�x�e"O��`��@n��b�35k"8؆"O��:a�T_��0b�@�-"Jt��"O��1c��-*��݉!�'K�=˰"O�i$��&�$c���TD^�Y�"O�G�9��e�Ս	�S�.I#�"O���'��Zi�����I��"O�Y R"@�3���V`�m���T"O�`�y��f�?E�D*��;D���SEC�v�:!�`��fT^mZ�/D�8��M��v���0� D�W�]zqC.D��c��L8�A��,�n�Pg+D�d@��D�v�떏[9c<�ە�)D���rDF%4 ��4ChZq�#D��#WC�Y�|�[��A�%B��T�$D�*p������)��G�̸�1�-D��CL��z�t�J���� %��G0D���/�W]xr�c�'L'T��6K!D��#�EO+#�dh��C�4�mjs�<D��BV��e�d\E�
��v�/D�|�@��R���H��9@��U�s�?D�|�`�_�+X����xɊ1���;D�lb��G<�ca�Cŀik�-D�xP���;T6ЀW:rW�(�"�,D��c7+=8�EA�A�FyX��7D�l�����!�`��z'��ce` D��ZEiрs��C��A:���u�3D�
!��4	 0���O���Vn6D�h!�O�#i�y�T�T�i�p-	�*O�y�W�Om�~���"��G?�Y�"O:�1�D�{ 0�bR��"OB�a/��Br�y	�3X�=+�"O�����R�.���Y���:W��p�*Oj!I�'�m����3Ƃ�����'��h+v��?��e��TVm*̨�'��DcuC�}m�=Ѱl_�N��	b�'ڭ��	��3;hA���K���'�D��͚{�x�{��Ɋ..����'�Хӧ, L�d܈��<x����
�'��а��S���Pc^(q���'�~�p�*��r-�I��A��ܩ
�'��%ڡ�M!7���@��M�%�J Q�'4�#c��:P�t`��Z���H�'�nQ���x׺0���ݤ]��4�	�'B�MrB+��,��.�,lY��'�B��� �$)�`+�6���*�'qf�(c��<��p�4m��� ��� ^$��%�({>eAc��k{~B�"O��Y��N�K{����n�^&	A "O�����5��I�L�tAH���'����2��\����D0Th�Y��',����H�.�(ׂ G�&�j�'�LX���04���J%k#@Z�؊
�'sR�"K8:q�!�sŋ��tL��'R6�!��Ul'���nX�9��iy�'�]�B	��A8ӯ׶S��(�-�/۪��R4�O^Ȉ�LK�R�̀ dʅB��#"O:IHd�ЙT�fR�̠,�F[`"O^*��/�y�GbM�a�j�T"O�|��-#��ˑ��u�I��"OI��KC���Qc(�;=���f"O��׭�:
b��AS�
�*�"OH�
�"��C�28��fۈ<���2"O�pJb*�+a��$	a� �"�l,�"O~LINf�xl!!C�J~ܼz'"O�h�k�&|���`��j��"O�%jP��T0:IB���c�d"O���ANP�u�Te��!�	ef��b�"O&,I1-�;������-vb�R"OB��FME�c�h�2`��,;r�{�"ÖA׬�/�&���A�-��"O��kQ�շEO���_:LF͹A"OF�J$�[!}d�`�D+DM1f\�v"O*(�4jԙx@���0�D�q"O>i��ܫA����P��L�"Ot1�u�Do�LxsH�����#g"O���0iH�^����ƅ��p�"O�$J4�[�@H�RVe�
Vp�Q�G"O�բ�O<,"%뗍�&�PIr�"OX������d)��F�X�R���"O���dG+6d�F1��"O$8��iD�
#6���C[2�x��"OtT�0H<S"�k�F~��aS�"O��
Te1P�<����(���2"O���B�&n�LK#�"b�J��2"O���L|��!I�$�  ���1�"O���шR�/tH��dR#�XH�3"O°�@���a���� +����"O�'�\�C�lQ� 9k�<D�"O��{Yr����L��r2�<"q����y����0�kJ8�&<+ǄB
$�)��6:^Հ�$�.`�"�j�@��;V��ȓ	��@2H�:/ؚ 0���M͘m�ȓv���T!. ���q��2����bʐ����fܕ�O�n��ȓa(��Z���;_Z�(�i_�W�x�ȓdB�S�U-����)p�����1��y�7M�>?;��(����h��ȓ(>(�!��9`������S�Q��{��$��Tk��)2�KM�܉�ȓXS���0B����5 �j[-/�l��� ����E�fm�e�d��0��8� k`���\���g֛G�b���j%�	p��&1�t��'�ZM��Z�� � (ڱ]
��I���.����o0��R��X����w���0�j���7�R!��i��Lw����5��'LN%�Q�Z%�v�8%⋝��̆���0���J �*l����?�zM���D�����
itѱ��ܾ��ȓ�h�q�Xo(�ȁ�J�O��`��S�? 
ػ A�T����%3|�� "O��p5��!d�V�1 �L��U"O��A�HN�w���Ǌ�\A�@b�"O*�G���9��!H�C:?1�"Ol��6jL�!c��Ц�w5�q�E"O����Ю|x(��� 'J$lP�"ON�sТi��Y�`��0ԛ�"O|��+�Ԟ<��n �l<�R"O�|�d	�޹r��)^�D�"Ob���Tx�$�C�y]v�; "O:����8b�̡c�#�9�"O����A6	B��+��u ��"O��
��#�����R�]���JA"O����#����e*Ï*�����"O���#w�N%C��Q��ء#"O��*c熅0��� �A˩*� j�"O**6OX"e;��i" ټn�H9S"O�(��ׯ�,�g�W�)J�I"O�XA1KOu��˖�-���+�"O�ْ�$�(!�+>w��]�5"O�L(�e#�����C�a��Q�@"O����)U3yÎѢc+ g����p"O��7�Ŵ9����̝z��0y�'������{�p1��JM&H�>���'�h�IG #��+D�./�>��'B�=K� ��@֪�냂K?��[�'� �b׌�}U d���cj<��'2�4���ƫ%���ڣ[�EX!��'�����K�MG�	�sɈ�;���:�'FH ��C��H8h�)\�4eD�1�'��d��l�
�d�R�"�%`��y��'��d��Q�%���m�'��Dh��;=��y���ߊ��'4�yI�eP�A�
L  �;q���0	�'�6 �G�) D�\�g� �YN���'�����ޏY!���%T*
4J�'@t5[BM�6-� �6�̬����'4��q�a�{���%�ZB�2��'(�(2�h��UA\�(f
�&5���i�'8N@J��҃P�N�V�
�*@&���'7�b��]HC�l	�H-D�U��'� l�q �"16��!�W5#C�<�' ��"ՠLna��˒��=ie6�Y�'ƨx��ጣ}M*��!&P�Z�4���'�Z�K�� F�����U�BJ�'��]0R�U� ��$�S5�*�''��0q��[�*�����	@�v���'O���`C�.>۰��"H�4;Uȱ�
�'���ۣ-��Y�dб�ߪ9�jdJ
�'��y�#SƖ�bQ(т,��@�	�'���@�C�B�+Ꮦ�%#���'N�`�ń�c�X̀5dH�sjFĠ�'�����kWv��w"ؾf
���'vЖ.;���Qce�>#XX����V�<�`�V,[��|��J�,�	�E�W�<I3�ˎY=Jb���2 55	y�<��H�/
�<��I/v�jf� k�<9�L�q~�dZ���?|htk"�Qe�<��݆Eu��X�M:���F��H�<�ID�\S%%7M)x���z�<�,�3P�Ұ3�L�2c}ّc�o�<IG�_�B��C��I/Y��;g&j�<�H�S&h-�$ުB9"EC���Q�<)�`��8`T�(s��v�HQ��CJ�<� ܠ�Ǣ�"5Z|�C��kD�ebv"O.}�����8�e�Lݪc:�d"OPi�)��̱#�M�[���"O�Y�
�fZX�P-B:e�@I�"OՓMC���;'�ކ����"O�� a�׍=��ĭ��TzL�"O��ĭyj�0a�>F��]�"OZ�A�NܤkI(��VJP�Z���sf"O`QK����e�` :���O��� �"OPmxrb�$��q6(ٳ^ ,���"OxP��ƃG�ʭ9���i��U[�"O�1�
��Y1|u �WC;���e"O608��G�f����d	5��3�"O�)"'@֜6Ix�s�c!	$�aC"O2��i��g�I�#��V�g"O�U�a�}�P�1aÖ�=ۢ�rT"Or�äoӱ}F�Ѱ;q7���""O�!�w�9T6�)AE[9��qC"O�q�rO��&窱�T튆����"O��ɓa�(7��e�cm
)n�&}��"O�=!vNC\����9l�%[3"O\)Mٗh����Gb�&Z_��c"O��C���f#���!��RR̬��"OZ�P�&�<W�m��b8���(�"O� M��j���p��r1,�K4"OJ�)��!KN�����(�"O���Ň&
�k�b"�a��"Od���(Ù`됐�� Q}4!��"O�����\�'�ڕ
���;�
q�0"O��'��>�091da�Ď�Ӏ"OxŊP'���d����+�p J�"O�)�R��0*�8���ݲ���"O�=	!C�Tj�3��, u�,��"O.a��f�<� �Z�'�8Y��0"OTU'f�9ԶX�fFQ?<M��)s"O��"׈"W�\�l��
�R͸�"OP �Q��Zv�Y�ڬY�P`"O}9�jĒ|��q�iFW"N�S�"O�����>_k 0 )�=���RC"O�b�	T�+~��"g�\��"O���eA�)|�H�g{Ra��"O�x��o�D�}�D��2�Ӕ"O`��iF�p�0� !��:�6=��"O4��c��Uf�a���V����zG"O8ܸsB��1n
��rmP�p�9D�#�E�̬�R��3�6�x��8D���f�/�v����b�t��A7D�4�f���څ)��#��x�6D� �Έhz�0���!�|�PC��+(wB�>Hrq�F�J��C�I�����b���R�	�7�y
S�:D�8��M�Kp�����jY��kc�6D��Q����{1�3���lel	���6D������'N���![+�Q��A9D�@#��/e��Y��D!0��sm#D��T�ǡP��A1*� j�	�D�?D�T��B�D*2�j��S�gMn��E;D�p���؄c���k��_K��!���7D���B�#�4��Aj6?!���*2D�,��Y�����(	� �)�C0D�$J����cZ����Cxt��Q�/D�dP�H�V��pI�Ɓ�D=ؚRg.D�؋R'��v��9)��}����(8D��1���,awn�����!Ehv*�� D�� �(�CH��FX��Q3�W IJ�"O��c�@�?}/dT�Ņ؀Hy��"O@D�w�º3֚�������"O��e�W?HĠ2S��$,��1�@"OU; 
�\�JJ�"7g��"O����+",\䧗�z7<�"�"Oj����.�ƀ�$��4���A�<�oǸu�4;���SUx�D�<����,K�u�.OJ����l
u�<1Ӥ@�F/��brG�,��h���y�<�� (p�z 	)<prm�Cx�<a7��8R#ء�&�ʯ7�,���COi�<	�f�tʬ��B(ܑ+��-��d�<��e� 
  ��   �  V  !  �$  W.  H8  F   T  �a  �o  �{  ҇  ޒ  ��  `�  ��  !�  ^�  v�  ��  ��  +�  k�  ��  �  \�  ��  � F � ; � �% ?, �2 �8 
? NE �K AR �X _ �e tl t " %� i� �� �� � +� o� ¹ 1�  `� u�	����ZvIC�'ln\�0"Jz+����K*ac�'b��2"��|:��MǟH��iѼ�Nx0͇I���F�
8��A���a������1$pM+�e��?`	B�?����挢SZl#��ׄL���>V9H׃�?����	r�@A��T2*f,��	@0�S�,��B�t$6�:��̆G��Q�#&L9*�jO��?�0�úI�<	zf��=���hPF��?Y��?����?�o��$X���L٣�`����?����?!�䙎�y��T>�yR��������cjeٲi��i]�b6y(�Q��?�����H�b��2@�C�U��x�V��t?���<9 IP1Ϊ��C�9	�)b�y�(P��.kN�DD����b�6FE��`�"Ȁ�Z�K��N�x���k���~��İ���
M�-y)O�rB�F�
" �c�֟e#,a�-T�3�B�'���'����'2bZ>a���X�~��A�XJ�r�a��	�0��	��M+��iz6�����ɿ��uA۴?�6l�b�$�7S0���cI�-�&��i��rmGz�K۩�?�(�޿:�V�Vd �ʤ��	�N��qR���8��²���%��a M�{�B`R�Cú��g�b�� �U� wp����P_���x�N��J����3Ud��'+�5w���
=f8��ѿ`�=Q@17���AԮl8�%C2�R�Ac�VJ� ��ף�l�	��M���p��t�xI�W,x:�c+�4Ajp0㲶���J�1)<��2�ŭBW��)5%��Qr"E�B����n����)��um�(q�/S�Q*�irl�M�L8���1nG\�A3a��V�JcßZ���I��ڰ�VxF�D�[�$  )����HE���A��S��i���%��I:1' ;IHNV��j�����7b����@ʓ>�V���0����_q���$�O: #1a�\��ISF�ܭ2EH�á�<y�C�;r�ı�OL��'� 4����:�`��p�CΓ;<pNa3�'M�(�C�غ@��'�. �wHS&U_fd��"-_~|�ÓA�������'ܐQ�I�4&�n@�C� b�"��?�����(�L�A�Κ%+�밨�>PZ썋���K���	Z�U��A/�=<�+���-byh��g��O �Ыn���O��1���mԲf�6���!Rތ��|�bO�.R�sǓk�4������9�<��ժ5�=��!�����������%�ЀY��!$��D{��DMŮ�B�ч�*:�"�l#�yB+O )B %��Z8�-Pf$�.�(OX�'ʣ<�p��Q��h�T��8I�	��Ƒ�Bz���3批tJ�#|�'�"��e�&�O��l}�WnX!]G�e�ҋ�L(<�����r�V0���ʐc�\�҂X�<)�霷)l �`�B�<��tjM]��p=т`�#'[fػ�i�"Y0|r!a�<�ѥI o�l��Cs��A2f�^�R��e�����{��96"���aFD�I�IA�?��#V�D娜�<9�I�DM���<Q0��-`��m�2sOR�{tL�7�yr�̻ʮqaA όe�� ��e��x�B�@����B�9J��%͞6`��B�IQ�z��c닼i����!1�^����y�R&�yBT����r��3Kh��=!���Z�[�t�C�O���"Q�i�4\�� �a+�f2���O:�Ҧ!�	p���$�O�A�%�F�QB����P ��4*����/�8e	�Y��xn�[�>���N�2K0*�aC��w��y��I�K�xM��� �f���K<0���'��6�O��Y�^�$+������=aHhQ�M�<A�������%?�p�ե�$8�GA�Cr�p�B�lܓM����'�	���:;�T$PcC��~���8��6_�hsL��P7^��I]�S�`���̓)UyP0�O�qzh�;�(�w����'�\�=:�zD�O������I�	� )#B�:sX�\�.�X��T�v��eK2�)�'#����CG#/��hF�@Yt�I�'GZ�H���?I~ʉ�d��L���K����bDǔ�䓐?Y
ӓDC�H��X@���
��;��eFy��~���3�,� u�Uh�^�N\��.P($����ˣ.zXu�-O���N�s�D���5�D6�@��h@�՗j�j��#M����A��ɏeD�3+�	�L��K-j��b�P���)LO�4�Wo�*'X�3����e������'���%�`��&��Ohʓv.��14LT�p�Qa���$�fI��'���c�@�2�m����F��%�2���<Q֌���r`�'��I����F"�5Q�y���0$�	
�xZ@�	ԟ���՟\��� �!kZu�I���D-H"�nl��GW�	
� ��V�RN�AK?;<�1����������0���Hqv!���@d���ȇ�φ]���waә<N�dI���N�~й6�I�:ۜK�i�qPN �0G�3y,�]�p��O��oZ̟��	����I���	̟x�Ox��G�X���� af�� P-O�}���i�Qh�{B�Ăiu.�
�^q&X:�.)���'�.��'>哉W�lxr��Γy�re�smʙs$1��${V<��'Ҭ��(G���\?���f�� �Y�bn� �jϗG����'/��
����T�j�z"�{��U8s�>
�ax"�T��y�|��7L���jT�Ły��e9����y�eD:.��M@N�F��
Cʇ���'�t#=�O�FQ���A)ז�!��r��tdG�S��'`�QYgD���yB�'��=p���6/�I�2I�+L������=� d������f-ќ�x$bt�����?Qp�xBf�L/48��-�^��!�0����Nv�	5O:W������pB�r���(�,��E�/����x�h�D�O��l�ПpF��m�I��Yt�.:�ᰂ�A�䓹?9���(?� 
�#-)ư�D��KX��PW*JS�'�N�I�'���	b�#iے��R�ڎz�]�w�#d,�q�VNJ͟4���4�CI�=�d���џ��Iǟ�9��
PrQ6'����O�y%"�a%k.}��Q�0=��
T�!�K�>�,=z��p��ꩇ�I
�@lr�g1�D�Afϐ�xO���O��DU�d�z�$5�<��*b�+�"�W��	5j^�P�<���'�������z2vp�S���J9��ɿGR�DA�L����{|r[�pX��G�nu E0��=h90���s�6<�'Cǟ8�I���e�E�U���ϧZ���2�I��4%
����2d����(Y��1p%<�O�As7�U� ɐ���+�`�D��3�������#�p>ن���X�H�k¨C�� ���
ڤB��a�����	�T�'���d��v��� �� ��&g���&����E�W���y�ǛZ��y2Wa�$9/T�'��� n���'P�rVÀz���',�pk𬏕u�	d��)C������'��(Z����'O�ƈBd؀0��C�t��	7(��1�'_}�����'������P��� R� �=
��ɬUU˳�N(|�Q[u�<�T���HB�z�4�oʟ�D�ߙ0IƵ;��\x&Eh�h�jy2�'x�OQ>Q�E��#զ́����y�8@!�3�Ɉ�HO�әU���@�4uM�]+!ʙ*}x8f�ןl�'����X�]�'��=$�8E�I7!����e����n�ġ� `Rh����Ȋ<'�(��%}�'Ku�'�f��ьQ?16�"D� �,��O��A.2�)§6���a��3� 2�T�\T�'?d���4'��e����8§?t��۲.Z*b��������$�,�	D����N� �4�D� �*A��� �8�S���*���c [�����cD!+�<��D��1n��	ٟ��	�6c�]��CٟL�I��0�ɻ������_��0���BWp�zDGПE���'��Xs��@)��Q��1O� ��L�Y�2��B+�P��!�"&I�	lt�5#�!,�3�IH��Q��A]�R�[�L~k,Pl���M����Lb������O�E���,g� �`EM�z3v��R!&D����#56�P�3 �uA<L�Tf	t�ߊz]�X��E�T�'��d�ҫ^�_Wl1h`�GPPf�1�,ˬ; ���'\��'���_0wWL�2�'�I�6�(X���	yb����#C�2�`Y9���`�TX���\��w�M x��R��ܓ2���C�E�A�x�k��7�O��`k�S��4�K3@1�� _����'�2�'�Iɟ��?Y��Z�FT����N
(�b���7�p=�w�� q���1W�ܼ1�H��o��'$�X"��'��'6��(7���������P���I=>GbQ:֥P���څ7�����Z<�q�4������;�X�IЇB.���"O6EK����t�����&S�9$y�g"O8�@D��uR)�E�ۛ�h�	%"O\ջ����u��IE�=۲��`��NO���iV��9�/�_XH<c4�6g�8,��$$>,��<���X���֐\�$y��	�B�@��G�t�ɇD��Ɖ�B8�|�7���R�d)^�;�Pi�B6D�d���+(|�9��o+�ֈ�B2��*�S�.Ö��� gvp����U/P��ȓ\���ׄ!/=�Y���1L@��Dyҕ��Gy�L�K(:�e. 5�}��i� ʒpAsM�N̓UBMD�t�e�����0@d���!�!3�>��#�"�PxB��a'U5	���A��6Ne�ȓVzl�����Jd�'�[5IZ�u�>�דF-l�����,��$KP�ܨsS`���˰ѫG��?�
��Ʈp���o�>! �	<��'����"�p�^2��W+N���j�� �U�0J^�2pP����H�G�T� ��2��
��t�P]	��� �,�1��Sb��S�R</֜�sDO ���N*�E	�&�ƹ�B�r�<�w`L�}�*%��Q<�JH��NR���:�{�J�>p��(e�cw̤��V�2�Ɂ�HO� j���n?��n�!yE$Hjc.�0�8��Wby�%�:"��<!�yJX��OՒ� w-D' ��*��P{L|"�'�$�a-߄g� 0�X�T��C��(O���@@8)� n\�#=�M)�	��y�E�>+z ��EM�5V���N܁��'Z�#=�OB(XI�(��2�ڈ��L�&]�2M�Un�L�'x5�V�'�I�c����.e�8m�G�Pe?�|
�DbD�O,IPP�,�x�A�;U�}q�;�H���*T��yB)V�?/�=��A�%_�h��PN����hO��̨��S5vg�m"�m-�I��"On�0���p����;
�)c�I�����}�'F�uʘ�<oR�����n$�Kv���$XrT�<�	�s�O��E�aK) +�\�1��F�(�z5l��.Y:�'��th@EÓ;nB@:�+�o��@
�'���6#^#pݶl�#�,	b����'ˈ�{��͈a
����u�P���'��,��
�/zȸs%�F�:���W+TA}rO3�2�qOe�1���z�~4��A�\a�(���'���BU����'$&�iQF��ߘ'�F��"�
�g�r\	��q�T�kC"Oܱ����6MB��;*�=YO0�H��@�0� x�\ BT�`�-m�<A�^ ��-{�a�MMʵ�d�k����{�֫TԒ�"Ff���<�"Bd�2��'hj"=��d�.B5�$�bLx��A�	)���a�����9�`�h?�5�>�#�W��@��D�2jp�Q�5D�� P��I������2sP��R�6,OԢ<Y�H�)t��ԧ��P{��C
m�<qf�"s�� ��%C�)±��B�쑞�'O�v��7m'0���g�+��F  ���E:��D�,I�I�!o=j��Ɗ�,�$�1%[> ��'m
��2E��p<)�UNUc �jf���g�x�<��-i��02��r���S��I�m���Owp+��Q�b�u���{r�X��'M�0æk�#\"-�2�<G�n=���DU}��=ʓ/�Ȱ��T�Lw~yV'�/޵���� ��b�ȋ�A&§d8D�`�G�,nl�QG�3
Tb�,�R���ɡk��r����5̊D(ء����a��6�$�jG5KIb��>a�5��h�5��m����+���*m��H��ɁEO�X7"@���P�v�@ŃD��>�$�ɍ��'�u���؜N���3a�>L�{�(�
���s̓x��Ts�D̓j�|�HF�\��xS�t�H*�'�^�BF��ZҸ�GM2^�*�`�'�Py)Wb��+9@�W�
�DI*6�'D��kV���W~���.D�"(����/'\O�y�=y�&5n����N��Wv�~I���QQ�A��~����~�P�sT�V�`|EA�fE�����7'J����ο>~q��£�d���
��ԻdP0I0�"O���U���Q"d��$h��'WQ�l��d�'p4v�[��
x(�DHs=D��;$�w�2��f�8��dY�);�HO�#�(5)!�>�F�Q�(1�t��V�.	���Ҏy�
K&��tj�#J�P���xծ=Sdn����_�1P4oMB8�p�`��9/|ޕr�nS�i��p���5D�(���d��
w�Q�S��0 ��2�D8�S�' ����&��iB>1j	יc��i�ȓJ"�`�4'}����GY.|d��Ey�F�>��I�Yx������/e�|�����N���"� �'�1OHP� �bnV��F'Q� � y�w�C�[��Q�R)�h�BቝGPU��(��y�͒���C�)� �r���	b,u`Ea� b��3r��,\OzL�Ƨ-�tcc��,
���0`"O�\�g�N��p*���Vu�E	3�&��D_�'� ���)�?{c� �A@#��s@�OV�hǧѿ.�1O�˕�Q#vO1O���1#\�Y���'	��V9�@)�%-D�@�GBO����ђ�(4��6�)$� �S��R��� d�ΰ@VوɃ�y�cI�p�����&�9B5q#dS��p=ɋ}R���BO�+����,���'7("=�d!������J<��ڤS�V�x��:$���!X1��K�1�IhN��>��^t�R�x`�54\ *ӄ5T��ЂK
����*�5Hn���'�Q�0I4"kI���oQ.�d�'b$D���#V�t>�S���1�<�롈"� �HO��#M��403�̫1I���ƴyb��ʐ�	%E�.�ˌy�#�3����F�R�����[#�E[wKG���+�$9Z���O8��	4GÒth�([�Cǎ��혃H:D��@�^T<B]Rg'�;H��b�=��5�S�'M�lX0ₘ}S��4�.M��i�ȓ#��R��w�j���M��DybN�>A��	DT���	\�+�^�H���*����J� `1O�M�e�ӍEs����k)]�Hm�Q]%1���)�J�v��B�	�K�����Wή�S *!]0C��M��5�AMM�Bݢrᆹ���4�I}��|HbߛR� ����T0�	�f&D���d��=5L�Gl�(X1$!z�kŋXo����HO���=��L~ʩ�*0�b�*��ޟ`��E���b����eQ%[7�b����]9�؁�Aɰg#��˂�
S�<y�ˁ�`��uď*U�p(��ʟOH<�#"��2�%�&��\��Q6!���3�x�0��j��5����4�z��?��Z����ŝ�R3���R)�D�#���:5Z�=�Xq^hcw�	�~)�va�%F�� �'�2S��)��'*�I �����:D�����֓c��,�4 ,�yr#��*BT� �ȯ^p��B��K���<���$_(W�(��-���
C�� !򤙛p��,��lj�����qO��FzʟɹUJ�#c�H�!�L��̕<�(Oˠ�R\�Y�x4�'�B�h���^�d���|(@�'�Xc������ V�DZPǌ�� �XD���m�!��X�O��ab�F�4%�4�F��>#v�'rўb?m� 	ϕaY4E�C���*9&��fL.D��	�*T4Az�8Z"dޮ{:�,��,ʓu��I:�(O"H� ���0�@%�F3]L,9�*9ߔ< �yR����s\c� �@�G�|��ѳ�_-!i<��ċf(<�̋<����^�D��3̚G�<�rOX�8�r�YA�W\�Z,&�~쓇p=��'X��qLՏ�`��5ȍP�<��	���`�b&F�nM�܊&���D�H/����{�"�itN� g�D�'��!�"�#�?a���I���<��(ʣ����<�&+�6t��GG@
�F��PR�'>PDxd^�t�J�0�)S�^�v�;�'�^a��g�f��A�0�
!N�b��:D�䱀�77���P�
�}\.�ⷍ:\O���=IC�O$,����n��>�zt�e��n�be��� .H�~"c��U�z��A������W�����$؁Ur�X��M�W�q��|���� �xDc��˭RVt#C"O��&	G>/�yYa-ЩqQ�8a��'Q�����9VD@���X� �@r��#D���pjU ��ֿ@_�9x��-�ɠ�HO��/#��WnQ���鏁k�j-B#�	F��t2�y������ X�<�(@,�jG�(hWF����xxΡk'��k8�\����@��"G��1@������2D�8*6N�8P?l� D A������,�$7�S�g�? R)[�C�e;��y��C�+J����"O��J�Ɵ�#����û5����I����h�'-��A瀙
�2�H&�&T������fT�<�r#\e�Oj:K��P8%F� #�*�L
�1�$E)6�ލ�
�'��4��"��L���"0m�{�'�0�FéD��1��<��I!�}��'��ء5e�P8nᨗ�ҷ0u��i�'p�dZjU�W`e0WL S�H{�]}�.2�GzqOYY��F�i	�h�0�3Rg�07�'ܤ�2a/V9��'ʊ�;cOZ���'�8!0�H�2t�T`�D�N /��=� "O
<q�D�.N�P(�i��{�����O�(1 *�s�6) @f՞m�j�QP�<���k�Qbf��2&�ܙ3��O��d[�{˗-A+½p�`��_(��!0c��'��#=�`d3b�������J�صO�ih@ ֐x>�	�q�Mj"� ��+���>�����08��xa���T��)��J D�(I�E(w�衣�10� %{&�+,Oآ<�QH�$DU���@�q<d*��y�<9q�E Y"���Fg���itB�tܓ>R���'7��j��ػL�4�pjG.j��B��,�c6%�`�D]=W�I�9��¤�^D]�,�?rJ�'!䙈,Y�p<����q<�sGJ�>E�PM�E� N�<Y��V�G��raJM72�P���,I�I@���Os�Af�<P����aJ�^�0	�'Q��K�7>ZH
?Y��h��I}�<ʓ>�T-
Q��6�n$ �i�|��D�#ho*Nc�09�h?ʧ�-J2,��u^�ظ3�B4!.x	��W*B�I�Z��q�ڶl�H�Q�?8JC�I��!2��U�3�vXa��8��b����	�L�@�"��G�[���%�B�	�^	� ��fOc���f�س	����2Q������XD̓*kz0�gc�yԂ�z`g�шm*F�ilxI�@��MT-
`v�$��`�����i���I��`�iƱ2^|�IL��\EƗԟ�i�g�zغ������ �H�n�Qx�V�5}��0)�(�:��E���N�uj  #��j5Xᣓ�g������+o}�h��ԍD����5̛&׈Ol鸕�'q��)I�J��A �C�Y�w��?��@����I���A&M@�z�bDl-}*�S�$��9�~¬B�%�[��,�{��ύo����'�N����"6��'��ӍI{���ޟ��nG�|���@D;}�0i����ԟ�K5fA<+0���D�}�HK�?a��;XY,�O��m��n��'�:�gM�����'��0�lΐG��haM�9�P�E��*�#n����ǲq��`�G%��y���<�������䟟�q�a,��G�TD�~��$+D��@����h���0���Zц+�	�y2���O�d S�{��9&M�*v�.��>{���O����6RP�%`�O�D�O��~�L�nS9`��7���2,�E�ѩ5�%b�	O"�AB	)m��[��>Fx2�ղ&/Pm��A�	��Ur@I�8V����Ę�XO�4���W�0��Ο�t���O�e�V�{"���,Q:Q�*?!�p� �Iq�'��*S�0�M�S0���� �A���DɃ�tr'�ʢ
�F�!D�`x��=B�Gx��r�Z��!�#��*��Ca�b�h�瓄Q"b��'�ߟX�����~�*�I�����ϧyM�(³�	 O�t�@jC�a\�ћ�ս5�$��7��7�a{����j�:]9�oT5�~ѓUcט=����F/�a:��;lO���'Un�tH	�D�;G�W�A:@Z��'�ў�F|r�Ŭ?hز  F�)Q����kH�p<ٳ�	"hʐM�1MT�j���a�lD!k;�˓.�lx����9K����c$�y6���t>iR�H�:$KE4L4��s��Ĩ	�N˄g����A�'BNY�~$�R�nZ<hArL:�O�Ԥ]�@�"������A�j��R�7���2Vo��(WJ�д,�U��̗OpT�T�:`��D��b���hdӈ��N�'�"�'�1��\��g��V���ȐC�� !mR�Y�4���3v�P2�#4qB�8e��yL��'�8"=�O� ���'�$�+�kܰwo �B����(��3.O �`�MQ�>]����O��'#NBu��?))T�UC�q(uc�8G�T�a����?�5�:u�U`��,8���?u� �� X��O�<��Q�2�����G=LH8�'Eb�*sJy>�x7�>E�D�����,ܘ\&U�0L�<�y�o?�?���������� �+���r��F�����01�"O�I@� � ��Ѥ�>���D���<Y0BDp��b���V�XYpS�*9d��,�9_�FE�R�|���
R��y��RP�V�X�1AֈJ		-Tq	��t�!�$�1sw�����,~*���	�%!�D��H���d��ULj���'R�|2��>NTpY�4/l�M�H��PxR�r��ʚ�mz
�x��P6: xa��Y����"��d�A)�+,�6RCҐ+e��/4�*�jb���'��b-���'��cem�0�u�r��E�����F�!�â&�R�A�B�
<if��R�a��Op�1����	�n��ѡa�_�!���O��R�l�:]զY� �8N��xr�9��<���$K{\��ZA��x�P�O�$�<��'�3�������?�O=:�j��f�����߻a!l��d��1�2�?��6z�$�v����O�$+˖�శ�N	^.D�`NX(r��x���2�'~�Nq��n�n2���t&���hF|�OY����
G�X�e�l� C(�g����"O���JĂ ;Vb$�I�jH�V�>���~:��P~?q�k��68%B�M�kcjd�֠�Uy��'�F`#�T>��g�z?Yg$��M�D��"Z�4��\0�_O̓]��'�"����B��9Rɦɳk�-&�p��'R)e.l80C�:=��8цǌ���)",�>E�VT�Ԙ���z�1"���
*b�؅��5�F�^�5٤�t ����M˂�Ό_|.ҧ�9OH���i�z�C�([�6=^}bu��:Zb�'oZ7�y�Z1����M3�ϡ?���� D(偗�[$���	0�Jo�&$�$�h��$QX���DBF�i��1a�a@=k��%�>IR�i�����$m�OUoZa 8��� VR0��dبM��q@��O@� ��>����/&~"~"E�@�b�.@���Y8��Y�B���v��[��Dɦ�9O���G�>郾iF�$���S5sBL %L��T�J� T��<�{���EW��k���$�?P�%�� ��ঠ@޴Uhؑ���5}*���\�z	��O����7Jd3�nکL[jŘj	2}�8���c�O��ʄ��` %�ify�}��S�MX���W��r�t�*&`�ȟ��4�i�&\���n~ʟ󤕲�������ԏK�J��iQ!P"��J[���'@�Q���7|��a���%2�	�	�'��lB�@޵ ��4��^�*P�ش�?�.O���E�D�'@�\>MBp�a�8�aW��3�FH��H��M����䓰?����(�t��`�����Ä��΀j�x��)�S,b���RVm�:l.�:�l�S�B�!4����CJ ��V���ЫdEB�I�I&�i�RXJ���C>�:C�I�U͠�� 'N9TA:$YV���7� C��P2]��Q!cx�XKg*^���C䉙h^m(��Y�{X��a��Fa�C�=�|Se�[�$U01�QJP�_n�C��$D�J��P�l��'eH�h~C��V��`S��H�Q�'��s�bC�I�0��Ǭ����MrL�6Gv#?	��?����?i�S����AOK��pH �f�2���i7r�'�r�'���'XB�'�R�'9�BS��ɜ���,�%��|Ӓ�$�Oz���O����O�$�O���O ��G��iS6�AP�Ko��x�@@Xۦ��Iӟ0�Iȟd�	ǟ�Iğ��	��l����K.�@�\�	m&$�W̎��Mk��?���?����?����?���?Yq�E>m��1Y���hq�-	8oP��'���'��'P��'m��'�Rd�1i!|��I b�;QbE�Mn6��O����ON���O��d�OX��OD����K�P��ě'"���S�N�x�mZן��I�����㟬��ٟ��	���*�E  ��4R#��F�J���Mk��?I���?����?a��?���?�v�X �s��96HJSaE�>F�&�'t�'�',��'���'���X(k���⧪���f|�'oG�9�6��O^���O����O��O����OR���>F�lP�5-�ڒvCC�DbEar�z���O ���O��Ov���O��D�ONP�&�I�S[$=P�	C�&� �Hݦ���<��ş��IΟ���̟��	���h��ϓp"~�H�C��>��D���ܼ�MC�'XHE3ŇR-g5�	x�Ld���J�nlf<W$!y���=U�~��9��'���'9������;|�l����Df�4�+d��q�, �I韐a�E��?1�嘁 5��w���H"n֪w��)����Q�$@�s.�<=8���ʑ�?yUB»?�P��=+\��'���,|9f8�TKh��a��Q�C&��DJG�y�@a��O˓��^,
P�C�HJ�ǀ �ܠp/�2MȄ�H���4~b2�A�'RpTy�O��'��'��H��O�y8p*\p�*�[R L1[BҬ�So�	-t�\�'	@6���Nr��1���8nL�S��8���92�0���M7��3c��{��QV�����O���l�41� ���D9?�̉*S����qDO�{��������`:$� )��4j���'��义��i��U�A���!ROxlR����'K� S�_�l+���7h:�E�H�j���'V�6��u7�C�
p(I3F-�6��-
B&Y��HGy0O���7B�7rS����	N,>�(�A���;�Fh[GeV�~�N�fQ�hJV��b�����V�(�}��`��w���r�Θu�L�`�T����ß������?y� E��sӨ�#`A[�"�x$�$Kθ���zv��r��Qwn�<y�[�e���D�u�Tm��u�IL�Q'(<T�V�*W4$[j= �ƕJ�|8����?���?9����$�#/�@Z���O�Ij7)V�H^Y�q��UD(	���O^LoꟌ�։;?�U^����4qK�v)�6����7{^�Q�てT�J�
Z1|���A�'��2gb��)4�� ��xl�A�w'm�@�;K���^�"��Dkޞ2K����\]��� ոF��'���O[Tp���T�'
~("���=y~�!����wIX	���'�2�';�( W�W�0��I��M��	� ��_�&$���-.�p�P:im&��e���0�6��k�AoZ�?+B P�-.�@�Mj��	4J��O�d����� �, ѥ��5�n���'RG�<AB�'�NiY�J ,n��'R) &C�Mңn� n�D�^B��'���-k�,��TVy��'�����8ZR�J�m�lP�!��2X��;!S�\�O��D�O����O,��Ӈ��Ԯ[�V�.Q[�8	"�p��FɫM�K��N:-�����<	Yw|t��c_�4�7V�����D�l�r�م�J/�@E��)�?1�C~�H����?Y���?������pi ��4�͔_�v�q�IL =�pI��A�U��$�O�mm�П`�2�$?y�V���ڴ#
��A�e���l�8Ce�e��i�8�G��bKhԚSJ��B��9q�z����)|����B�$��`XR�E�"��Ր��s�uAp!���?���?��'-O�C˟j
2�ɮ|\�y�Q>��2҂-2:rMB��'�"�'�DeQ�����'��7�c�����D�
z@��� J�N�;a.@lڏi�,�	772,h15�?��q��t'��(��ωE��yX��FPb΀�! ��I�
|dHQ�'馜HcN�<	��'�Y�a�[�A��F�!m����F�=��<=���	ʟL���d�'ڤa������'�B�H�D@����K��5��2U�rI�
��\}r|�qm"p�
�I(V9b]cSHJ�֜��-ǃ%�
�2�K�d���D�'�.%��O��qB�0:O|�E�(���4]��{�d�����FB 2op���Z��?���?���ȸ���yN~Z���?��'��&���yFΦ2#��#�@
�k�ʄ��?1��=1�6�'ԨDi�O��iƟc�V��cW]���y��ܞB쾑�3@�|��mZ2�|�9���(?ǔ�(Bx��&�G><��.���'�&d�<xr�C*�0�Ӣ��!��$FϟЙ"@�q�������?���Eɔjfe���܉d<�Hb6Fƒb�'Љ#�a%	H�'�B�O%@�Q�T�,�Q��l�ha�a�B�8�ZA1��˼���ͦ���4)��T��wSV���D#� �T
o�m���nH=R�@	@�ָ�6���o�>P�1O��A�b�:�?�fB��e"�4�?���)"깉��\=X��{����&�k4Ņ?�?i���?����?�-Ot ǳi=�ɭvb�AY��� d8A� 5�إ�ɳ�M���xd�U�']�Xf�m�V���K>$S�k�o3�[A��v����v��V���8u4O0$"�����u�%զ*Jܥ�O�ݧ����	�p@�¬XT�@�fY`9��D�O���� ��37�	�O�A��Lʳ�- �g��E�P)�l�O����Op���5Jn��!=��'`���'!���p�[4\���*M4&� Cbp?�U��)\� �	�?��SM���z��U�a���'�]S����ƌ�*/�����>k&-9�'�V�HF�<���'�h�R�C]/]�B�'r���/d: r�CG�1��3'�"�'��ɴP��`���ɟ��������K���#c	�h�p�woF:��ѓ��Jџ���>�����������ð�ٖ'H��Oe��2SM����fVI��@�񈑨*�B�Q4I�,�p�͓�u�I��y2!B%��(&��=�'�ۢ\Fl#�K�)Vw�p����Ҙ�Ɍ�?��?����?	-OJ�3�W5I>�P/Q%+�&�{��\3
%��O ���������W���|
/On��S�0C�m�$* ��i���:@��7-֦fC���R�l�
|KE��O�(&dߋ�u��
~�%̓p:��@$`	���d��L�D�|Tbٴh�2G��	r�h��'��'��U$+����,��U2a�p$0���lO�:�t͠�fM��d�O����pHw0�&����%λe��dh�㙧3X�PuM� ���Q��M�dC?Y�dP>P����?��r�Ƚ І��F!M��2�l��8A$�[&�)fy�I x��S4O�M����<v�'�@q�"�B%
b	Ըu��+fE=�fC�Q-d���'A��'��I33d�ra���L�����k���rFL�B�C5�n��5����c/?�sX���47ɛf���~��%?���.�-|���P�;1@D5r�a��<�"�i�nD��(-�O��y��'0�p ��^������O@�*�J&8R<&B�O��$�O.�E��]#����$�O��	]� �CP�G7���@o	=�d�$�7jڐ�2��O �$�����	�bF����ӈ,e�Y��iC�C�7w�� ���cv�ٴ5l��ʰ&�:�2�O�<qsm�*n��}�����J�68�� �82%�x��'?F��'���>OGjX���O@���O�	L�ɢC!�,7���x�F>]����<�aD� ���?A����h���d/D���Y2J�=<�ָ!�S�F��)�':�7m�ۦysM�����,���	��@M�cn�<���W ��hc����̊R�D�#��7{��
�v���'���W�4��H��#���l��DQ�M�'zޔ3��6�D����?����?����ŖABe鲣g�� D��F�ʕz�N Kd���^\8}bs�'��6��OH��s�����O��n��M#6ꑨ6�R����0h��d���L�s�`k�+ҡy�$zǣ�3�?��K\0c�Z�]�+n�`:Olם��y��T�sXݺ�o�� .=ˑ�<��L2���?���?	��Y'fhkM~��s�������d�&��g��?a">�:���?��f���Y�
����dK��9���`I`�	`�,���;���H���:6>�`A�O�*ʘ�(�7�蟸��/ķ;lԠ� ��O� �Q�'aLY��D�3���� �#UmБZ�'���T�HJ�i�=SD��?9��?�O�]ԕ��,� l� �j"�?a���d"3I������O����O��Ɇ#4�X̂�I՗m?D%pV/�*z�~=�t��<��S�|�I۟���@����GP�8'����(�V���d^�e"$���)&�f!��m��sf
1��(�<L�$v݉H�C�O6`��ECRy���(N����\���fP�,Z`E ���O�ǧ�Q���D�On�d�O�d�<!$H��4\K7b ���Q� ��dH��a̛�?Q��g���'�2���^>�C�Ol`lZ��2��ۚt�̄��0��x�شM�����J�P
���?!$�;9�F�݇0��ĳ&9O��q�� [9p����[`lʠ�Ӱ)���>�&�`	����	��+x4��O�d��A��h.|�qg��v�ъ���K���?�����f ��|��h���0��0��kѧCS	����|�d���O7
�:���D�I��OI����\{�dZ��!F���ڀ�Q��|}h"#�)t�b���'-���W���<qg��>�����TKw��%�����K�$�"�%-�:�4���j�O�$�Ot�D�<�O�c 2E�-O���Q�}4hɐ��V�z>�)*fa�3d����rj�D�O�'j7�Φ[����@��� �fP4�q��&nx��`�U Ԙ#t�O�����TWn2�[LT�k��l����Cu��Z�P4�n��!E����heG�M�x����?��P+�(��*V����?����y�k�8��g���U�n�)t��8�?��"Q�e�J-O@ nZΟ�'':?���T�4��p���C�L%8��D��b{y�F9����)ΌU��!`���<q�C�2����7�n�B㠇�2�\@��HۈO-�PJ3n�![d�I�?94�]7)px����?�������԰�`� ԩ֬?gdH�f"4ڌ$q*O�iDl�<:����O��d��8���D�#0���5u�x�aJ�*����'�7��ЦE�6m��� eMX���&�(�qI�	�8��7��*l�Y��fَ�h"��~��:R�cr�޵"��i5B��^֦A�tB6ix�E��Ն	�#\#�uڴ�?a��?������O"-�$a����O$��&�:��!$�l�ձ��O�EmZ��p�I$?isV�lQ�4Pq��A�:Xm̠a�iX��s��ωqK���]w���sa��y�D�~�Đ��`xZ��FC�|>��8c	�2�4��2O�{�i1�G�-��d� �'#r�'��4�S�'��O�r��#]1 ���_g��("�!�"�'�"EݞI|��6�':2gӨ��]?
��$R�������1K~j�k�;��T�Ox�2��`.�6-�d)zԥ�1K�v�z�<O�#�M�fP���3�X�8%��B�@��L�֐K�'���Q��y�/�&�y�c�,�?��?Y��(����O �b�l�ib���?�-O�*���i���O��d������A��.�3�Ǝ�,C�]�cm���r<�П�mZ�pcJ�	�ZJp��aҟ�
����B���JڵI��Q�NC#@�@B�TV�4�)�'��Ώ���U�Q�˓@�lx�6��0}yT�idf�ܲ Q�'��8f攸xQB�'J�'y�W����V��C�5i�B�ַ9��xq$Mhy��~Ӫ��G�jL��"������Z�-}7
���l �V]� R�GR��M��Ϙ�{i*�!�K?X���X�����x�m�j�&~[�i\'��,
"N%if���v��K�O<����Lr���O��D㟎���f8�����F���(���G�� �ɥL�!���Ο��	ӟ���:^
���۟H[�4�ygB7,W� k��>W���)Q�7'���jӞ)C��Oؼ��xo���O�xH"JS"j:���E��@���s,�zSE��A�S^��=8�����R��-O��	n5�La#��ߟhr�1:l��(�F b���$�ן��I��	Tyb������6�'Q�'��S�� ����J9d�6�'��|��OV�'+�6-E��a2��P2�Sb\���@�
�H�
���~�h`��2O@�H�xU��)̔)R�ӓ3�,����l\9w�]�s>T� 3��"6���`�?�?	��?	3A�;�(I~:���?)�'۴�y���{|d`��ǖ��^Y!��̺q(��D[��q��`�����l�7v�j8#d��8"�tPY�	Ջl℀���*Bt�f$�ʤ�;��٠1=���'@��#�`S�cƨ(J�}!�	n����̅�9��X�C�<���'͒hJ�Z 3��'ab�O|(��tf\�o�l*Ă�{��PΖ�~*�ɇ"'����������矔�S k�f��'6�Q���<����F�1#�@�R���>I��?AjEi?1�aX�v \�'Qa���pg�t��D�OI~E�C'ߌ8v2u��A�<Q坻4u��dR�9�*��'����%a�K%"�S��⁶>�mI�#�|ɦ�d�O0��O��ĭ<Y�O��=Z�!��7��b���2+ļ�%gNXⵋ��<���'H`��'|̹>i��?�s`���#��/?NX�chƊT��u���Åqi�%�)�?�D�VA���݅BC�mɄ1O,ם���Μ��յ� ^�D��C�V�2�]"@��< �މ��ҟ�	�?M�vK���̳��(^J(�R�FXVHXA	�J����I�i����(��'3x6M�O����O�h(�I������z@����/�~RC��>��%�ip���/���զ'�yR���B� ��(�X�V�
��44�E��ΟL@D�^���D����RR�L�h���I���̓�aB�OC�����Eϥ!Lu�	�8�'����EI/W���'���O�
@��K�	��<s����x���1&��k��	&��D���}B�4fy����^J0��@�?u�A	�>)5|5� p�I��A�' �5� H��Pd�dj�Ku�Я��> �	�&�2��/O�Q�u��?,!Z<�IkDM4n🈘����P�d�������ß<�	[y"��)� ���M��-Y�}���3��(!��ܾZ���'�T7M�O��1����O2nZ%r��b�Z&�4��U�W
D���C�4_���u�@8�BE���?YӪ�@:d�]An��D7O��B�J�h$n	���/��̨�@lӦ��	�:,a� U֟$�I�p�S�q�L�O"�I:V��sr~7�R?�"���g@����F�'0b�'B�$�ňM��	��M[�w���r��Η:.���BO���и��M���z?��&8Jl�����?�	F�
��A2�!,K���'L)	ti�E�7y��9��>v���1�'@Bt{�ļ<���'� r����~���>H��ʓ+�	x+N�]��O����
�5�����O���=_�����rF��Pw�BJ��$׀Ig�ɡ��$���Q�ڴm5�	��8$B��S)�%S����l �3,�`�*�\�\�9x�8�%E�_�v�@�|��"�ԟ�"���Z�yQ Q�c��5y#�G,��@�1�|2�Q�����Ǔ{t�!9a�=gJ�=p��K�C����X��������	��M���H����'"��g�6_�d�zr&^ I[�(�ʙi��rG�O��7-�7����큮mz-��9O�d35���u���.�؀1fN��&b��"l��%"AsoKOyr(�OB���/M6 �����O��$������ѿtLX���jݽY�ƌ�򂓠�~�l�h���͗>�?����?��K��a�'�?Y`�G�ұ�6�R�R�P5�#�	��M#ѿi��x��'����n���Z��'�VX����z�Y���P�|�@!��:�H8�@��<)�������9m�E�'/l��D�R^����;���↓>�8)��	j���O��D�O�d�<�� +�!q��`�A�:yTP��_� ��)k�&��'S��#�'�l�>�!�iaz7�@�='�ɑ���0:%J��ңo:�����\V�9�� 6"�$�4)����^woD$��cb�$${�=�S�^ġ�%�	(.���mډ(Șc�d��X�V�)~��ݲr�q�� ��)!f ��O$�[I�H若��|j��i��%Ɯ�~�K�:�b(!`G]�~T+�bO�3�N���X\ ���V��M+����eXtGV0�a̓0�d�3p��|!n���IY���R�H",�����`H�[�����X����?���?�F��318D�d"P��B!�Iɣ�?!�����A.e�d�"��Oh�d�Oj���Vˈ,�6A�1M���*���YH4�`I�<�X��y�4I�����~"l"�ȱ�'(���B���S���4���,!b��vv|�Ԉ�y��}ϓ�u��^��?��O�5��	z��1�(<�b�Ҷ#ɨhlH��$����"�?����?9��?�/O������Ikub���$<�9�/ɘ(դ��ƫ�O������	����r��	��M+%AFh��$�&��[�XX`%�<���"(�^�jp��8����'ݔ��r��غ{1b	�t�	6c�����GM�|�J�υg#�<mZ��?��I�U������?Y���T�������%��y�M�X����!�P@��lB�� %���'��O2@���]� ��4�yg�&~� ��R�R49 IB9ԛƌb�0H ��O��Q�aw�4�O����cd�p��
�T�i2��$���E뤏^(d�b��'NV���I1{��ջ/O�P�I;h��3������(��4)��I׮a� ��L���	˟L��Eyr��s�
���'"�'���p��[�Z�kҧӀ4 �ZQ�'.Z-J�OL��'�^7m����$-����d�M�l�mj`�OP��AA[��������Odآ�	Έ�4�1�57���fݑAs��OF���$�ns���� Ľh��F��P����?��%�`������'�?a��y�j�>To<}z�'>x���E�X�?��d�@��/Olqn��|+��!?!���5��%Ru��ѴA)#1BaB� 5R+p��C��O:�j �r���W�l���Y�.�jIZwz�]2�W�8C41�w�P�N1����B͢eR�Ք'8���&E�0���O��D�O���(G�ڈؤ��Zq�,s�ī �,ʄ��<ɣ��_�]i���?��ҦD[�����6�*m�rƝ�m�*���H��Uߜ%�'NR�'��'��,
�[Y��+P8y�~�PV�@�j��={�j�H�L�����wh��b���S���tʓH�¨�	�A�T-��.��$I��2����C#�2�'�"�'��Y����A�#"~R��	�����qV�������I��MK�R�0X�'s:��?1�Z-8\���t�Ƭ �G�P|���,e+J�i��O�q�l�z�bb�:�d�$,<�a�1џw�D�aȆ.kP�#�-T�{����l���]���?9����#'����?���4&Ⱦ����/E�2i�u��	�?Q��?���D� �u�.O@\mZ�T����Ŋ�(�R\���7"�
�Q��ѭu�d2(R������
� A荅>��R!��OB��
ٍ!���,��3j�:RÌ,����*� ,1�T���� ^*�P�N-�?����?���T��U�q�Q$=��MR����?����$,e²���*�OF���O��IE R��0���dghJP"�!٬Y�!-�<��Z�X�Iʟ����`��PxW��Ofa #@Y�8����I�}Wd p�K	��ÄG�I�!X�4O@�]�$�:�$�a�,��'�D;�l��.Zd:��R�	�X(��O��Y�-O<�����O�D�OZ���<���8M��`{�å89.����T�Q��9!�N�*�?���&=�F�'X�+�O�-�'�6��	.P|z�g ��[�F��ƐlڛN?v��C�V����m�џ�x�h���U<� 4(�' �1��;3��j3@O��M��M���'��p�%��i���'���Oz-{f�?�0���a��Z��ޙ)ǖ���F�*>p)�i�O����O��)J>
��)�O�pnZԼ��oc���w
-���jW��M�w�i*�a��'�Q�k@��J��+o���Ǯ�
�$��� c�`��@�\.�$i0�6�?6
�GL�D�#"�LT�'��DɄ{���K���O�-����l�faR,�sHV����O2���O<�d�<Q��,�*�����?I�N��d��BK5f]�T���҇K�,i�F�`��'���?a��I/f��'�80�V�ă/0�%��O�8N�0��+!#z��ɲ9�Ti�� ����]J�Ϧ|���Cß��b�B�]���vk���D,�
�/m�1��'���'T�k&���l��O��'��� �͠ ���.5I���>���v�'��� �.lk�I��M��8���'��4��0x<��!`�>�Zu�.ۮ9�8��UNg,���<������߰&�he�'�z�������/|�@�i��ه}��c���+�Ă�Ƽ<A��'��CK�*QB�'���O���ڣ�H�W7
�p (�1q=l�k��	t��,L��]s �F�����Ο0�Ӕ�>��'�v�`��"j_Ʃ�$͐*G`���>���?�c?��%�^\��'D��m��F���ʈ��_�7 �MB�(Bl����T�<i�G��Dہ\�|��'�x���!N�p��@A8^��bdN 0mPPK�eJ�T����O��$�O��d�<!�Q�\����,�d�/�jmza.R�|o�����V�'�4m��O��'=67-�ۦ��g�
�G25��圈/m���r�i��B#B�u�H�avm|�X5��N�N�/�p�[.�t!�;p�(Q��/(H�'� P�kd��"/��A������	�?�"�ƚ�S˟,S�#%�����IY��$p��CƟ��	ϟ���� t��ݟ �4�?�gd��<���y;�1�7���GI��DI�/�]�)��h��K��M��'l��)�%�ڛ'�����|���k�#�'G�,Yzr�Q2��a�A�G=`�d�3�bT�'��$į~tp�@a�O&���OZ	)��X�C7x���OL�w�<@�3��O����<i�S�.�`E/O����
%�$jܻ`�T�+�F��:X�tC�_�+��4��'�M[Ǿi��m��'�<�@@��
Qₑh��ˏ'��=��Rw�!��g\-f��Hx����;����qBDt�*OY���X"��A@��Z�(�C��Eӟ��C�Ɓ�J����h����C7GHy�S����%��)<�hH44f�<K[B�'��6��Oj��Pd�|
4T����$Tj�su�=9���S׫D�uLDnZ�wPyj�D�"X8������̸PU�z{�H�F��۞'7�Ua�"=n� ى"�T5q�Ѐ���iT��(Pf%
0��Ot�D�Ol�i�9��D]��;��3(K~쀖)
,
(qCE#�	!x �'�R�O34�9��'9Fa����Z�@)�)�W��"�+%��æ��ڴ
���r}����?���8S���W��z���yë]�PΩ��'Y�>��A�,�ȟ���	,8s��j)�<9G�'�v���H��y�]Ge��'BN`'�d���;�2�'�'��	$���p��؟ �I�����eբ]g���o��Ah�a��@p��r��ɱ���ۦ�ܴ#�ؼ�O��@h3�U�Oɲ�A�L=I��I0���y�F�I b<����أsB ��0�|�$�[��4i�jV"D9D������ ��F8��D��'B��'�Դ8���]��O���'���M]�ِ��/jp�����
�=��f4k/�m�4�'���g���d?T���?�0�\�t�{%"^-�����V<	+@���ɪ�M˒%�[F$5`�����/"�)%mz�	� H�^)�)hf�B�|W�H��� p���Z�U�����Mު���F���?9���?��'MQ���~gv@QEm��$���WnF��$S�T���k��O~���OX��I!xS���O��0cF��o���D�T��X6�Dy��n�]c���rrU�̟��äŋ�rl��4��j��N�j����4&ªM��Γ]��MH��j�<����Zy�OR���eZ	f��+GO.;8vqcǕ)M0)�գ�O����O�d�'�M�&��ʓJ���3�fW1��sχ3���s��.�$q��	�?I�ir↏��y��' ��'��Bu������V�@:��2�F�a&؜zt����uXx))��O�Ih�A���u�Ds�����u.l�Eb�H�(� ����Q���nW�z-�Z�@��֟���!�r}&?�p3��5>� "��8��R��;9���	ϟ���!?҆��F�yyr�'������y���%<!�m����b��#��!!bȡ��'�����6��F�O�he�DîP#�'m�<��c�����z�o- u�D��C�&~`n���+�BD�.O��ɑ1_��*6Aןx�	ӟX�#�*kA~1����b�����ޟ��XyR
�
Hݙ�'ab�'L�4� \�b9�$+E$~��R�[.\��]��J�O\�n��M�a?��X�`4�S�_��s�[=$����'�����ۭ@��;"k�;$��dz��7�O�(�h�Ty��_=2H���Sұ{��V���d)[U�H�f��O��D�O����O�˓ ԰��B�(.M
5J����bʠY�*Oh9o�ԟȹ��!?1�_�H�ݴƐ,�EG��s_X��K�!�F�i���E$M8	��	;�M�y�߃YĶ���v��]�%��?e��ߕd���i֛r���%x����ɘU���B`�L���	����%�4$�O��\;!%J�N���T�]1�>�C.T;N�:�����?�����&��|��k���'��T9�iL�^�~�JK1w�����'�"�	�~2�T7$�i���B�N7#a��1R�NHN�rS�ئA�#�FS��s���46,�9�C�O an���d� ��O�����(l%��J%�"*�(!F"O���Eۯ�PA�_Sx��;OB���l@���q` �o�>�a�ę���dǷppQ��i^�]p��C4Vo\�S%b�! ��!�6pX6@X"oV^����b�x! �*j�u�d�;��J�	(�q:'�f0�`'�_ސ�z0�JMbg�څI�%nd��e0 �8� ����W̸$:�`Cgh�����3Kkr̨��ē�6��'�H�X��w�ʑ0o��hc� n5����'b:���b%�-��$��:��N���$��Z�c(f��@$C��t�0)M�e�ePf�G�g2ؒ�LL0��T�faYs
 d�Ǣ�"W�,a�*�V�2p{0��F�@��'��	 �:�ʦ��9�!���#O� ̠`-�b���:���j���R����jz&cDЙI�(F�Dl*�S��;Q\Ԕ9S&�^���g�;R�����O6�d�O�������Qv��m��t�E�i�1AVc�-��D�.R,r�'S| ���'x�'+�p,`����:X��|jVA^�hoW���УL��M����?Q����#_�����S��V�� ��25���X�+̌��@�	��0Ӗ)L��2C�7�$=S��gO7AN$��B���?I�#ϭ�?i���?���b,O���F�O.	��a�:=a�]��+ް	�o�OV\���ɬG>c�l�����U�Fn���i�v��O
��	�����矼;+�ey��H�)���'��)E� ��SgD�,#��{�j@�5�h�x��'�'?�\{E����'B�'qm���Eט� PɎ�k*�I8��'+���9\��ɚs����IΟX"(��杀@�H|x���|���!�F�z��ʓ4UBA�<����?����Vmw�uj��]+,a�X��E�N��vL�<�s�S��?1�q҄���?���ɟxz4k�<nF��Pt,T��q�	>f���'�������Ly2L�+��	ًWg�!��n�_�N��-O��"���y�'�b�Z�b���?�w��yB�*PLxq�q)ֽ|�rBe����O��D�O �D<�1�/�(���*?��@�5$ TJ�U�!�ɀTg��$�OBd{S�Opa��'����'&�1O0mÕ$��g˂5{q�\]9b ���'b�'��I	̨)�O���'^����BI�b�	
eϜ;�"�h*t0�'�v�p���?a DYw�'h�Xt>Df�n�D���T��RW����!����Iܟ��	�?}�'t&�Q��ݭe�&i�D��*(Q�(�2 ƱBnb�'f�<#U��&3��'f@�S� �2'��ե_����A^vT������I��$��My�"A���-L�L=#qbO�F�~q�K2.�j�("�Oڝ¡���OpYv�B���{al޷w@�ٓ�^����	ٟ��Ɉ�@ᰮO�(@�=OD�dÅOQ��P,�KP a�UD޳JJ�Bj"�I�(��I$����ԟ$�	"&dAq���E�8 U+��kD�4��ԟ�a����D���t�'��	�qW>E��JU^:�gE<62+����'�Җ|b�'��V��GJI���*���4D4~݋�N�Y���)OJ�W�'���[/����<ɱ��#k��0�I�f��EP���?������O��D�O�˓=�����Oa�93�N�}�<	!��em+��<!VeP����	�j>@��O�i>A�ɢK�=p@ �.�,��-J�P��0�'���'��P���Z5Qj����Oؙ"�(�҅U!t6����O���_O���k��i>�	���&ieaħ5:yB�(�.Uy��d�Ob��?��5��i�O��dc�Q�F�&.�2!7�!H�P��܊p��$�l��5O�Ԍ�(�Od� �O� ���葖\�F��o�<	�������?����?y����@\��RPq�9+��\*z�L����O*�	$g�2XZU�)�ԍX\MЅ�Cl�wh48���_+�?a���ަu��������?� .O�9Q�O�@��vHR�4u,T�@�]�;�6���'�����'��|ʟ���O�5�dBt��)X�Ρ����N�æ�������I% O��k(OH�)�O�o�7s'f!2�fE���a����(8�&,KA�'Cr�|�[>��?�'7&�c������JC�-)4�����?�����$
�ir�����O����$O� 7�@-HGZ�"���J��'��1وy��'��I��j�O��3��*%$�-+�_�ZU��'��T���'�d��~�'�?ɘ'�H�sׁ\�%���YB��R�A���D��'?!��?q����L^���=oT�j��O�K��#�̄���I�z�����O����A�|������O�pq���dǠ�* �W�=��d�G�<���?i)O��$���~�'�?y��EY'�D��
&��F��?��'oi������|��.����'5Yt<�s�3�B�ʢ�U?E���O���<�qj�/i�꟰���?����:��*���>w��*�(�{�f�	�r5����� � �b��&��̻Z��I[�[�h@�5o���.��	Zy���0�T6��O����O��HJ}��Ĝ&��\��a�7O�
(c���pw�'҉� �yB����'�|(KN?����t#���u�v�����O��K4�����	̟����?�Ovh�7O6�x�&�\��
�kΆB�8�����O\=����t�'�l]����'�����:;�]���
y&�,�aoӬ��O��d�*���'�>U�'�OU�MV���ӏ>5Xt���&NX8��QU�Д'�vE{�O�	�O����O���G	�. �B r��E�~3���g��O����H���'U``�'B�F��yB5�Љx�I�5�葄KE����9 [�����s���	쟐�	ן��	jy�L-D����.��� D�1,��qP-�>i+��<i�cۖ%����?)�#�.R�(�b���U��h��I�o�L�'���'���'A��==,�p��P
0����,2DbȾt�2���<�������.m�<�S֟��I����I�eRxy�&k
!I(A��j�tH1�	��D��៘�ICyR�q8�꧂?�� P�����G�-\T�J[�?y��S���̓@-(���?�v)��<��|rcƜ��5��e#z���E��?���?9*O|i�Qn���'2�O(�B�c�.���b��w�0�S����y�( ,�'Z�`�'��R��ͻ��YB�	�_��A��0�:���ey�,ެ.��6�O>���O��)X}rIֿ@�4Ye�	T�R����E\(�1�'QҫZ��y�'��I�O���O� iX�����q��jİRp8�
Z�B��iN��'B"�Op����͓Y�ؑ	 �ޝ+M��Q�F<����:�\�̓��d�O�����O|����<l�=[P�P�Vq���G�ۦ��I��	�{Qj�O�`P;O��$қL�t�0 L�C�:�A��M�3H 
��O���<�q�����'�?��?	��\3s�L�S�EHTH�(���?9��k�0ؘ�T��yg�l���	a/d�	߼�����%7��u$N�ܮKk�	\G��	쟤��ɟP��ܟĖ'���l�
�`���Զd2
��`�030���͓�?�S�<����?��̀ J�(2k�=O�<lP7!�� xH���yB_���	ן8&?��7�W��Ӥ^=��40�
YH������sƈc���5bI���?1�I��$h̳��`wn��;�d�H����5�2Py��'�b�'A��C�ru௟��D1{�� �o�}��t�p��(���D�O�"V0OX�)��OF�$|�qOL��B�W$Hل����$#Z�M{���?I*OH�rvY~�$�'�"�O0�$��L��e���[�����L!r���y��<r�"�'rD\`���d�Mx#U��,�6�1Tg����$�OP�$5Zhȴ�i��'��Oa��T�X��kEM�)��/�Z�T �W(��?��b�D͓��]=�褟JZCnL"�P�(��V�$X)��'.�H�eu�L�d�O����L��'���K�'�|,r@ɂ{�Y��Ƒ2Y�p�&�'@�a�'l"Y�\��%����i��w����5!� �蔎w7��O��$�O­ѐQ[}rgE �y�'���s�AкfAP�PZ�	�I[�q�~���'CR[�`��o�c��(�	� ��g�M�@�K�x�Ƹ�6M����	�4���OЙ�5O��䒢$��$}�5+7�)!P��nѳ7�T�P2L�O��ԧI��D�Of���O����OF˓[��ճ�hˊ$�6�X�?��1�f3G��I�c�X��t�V�s����ߟ���d03�M��(�e�R�T��@��/*?A��?	���?�(O|\�"�?��քǡ?�!W�B45��6l�Oh�9�7O���<U�������O>�C9Of�*�Y"X<t�T+ْB5�4�%�<9���?i���D�J�B �O���K����%Ϛ�J}ʔ�͡v���'I�U��'n��'|�O��y���ħB���iʌ�a����T-�'Az��'�rY��*�ʜ�ħ�?���Ed������7]�-X�$�[#eI
Hy?!f�����	�i.�Io�	ڼ�#���r��q�6Fm�Û̟��'<�}��g�R�'�?�'L<剄6�pF���=��d�4%Y'$�ԩ�G�OZ���s����.�����8r�pa�֘h���Q0�ݕ> ܭ�I�J:��4�?���?��'����󄆲l)��h�!V>T�~5�Rb)*����`�`��7��Y$�1����^,h~y�g;t�+�N	- PB�n�ȟ��I��lW����]�M�2�'Ɋ�4b�+�Bx!�eq�	1�&I&Ҙ|㈳Z'�Or�'����ku>� �j\���1a�F�'�4 q���<I�iݟ���?q%��:�ҍ`�jY�!�����k"�(O��+��$�O^���Oʓ<��:+ǿ!9�XYc�δ-ؐ�������Ɉr�����O<8��?�����<���_'�Z,Iu�\�q�l���K;D�f�	Sy��'��'M剕s�X��Kr��c�ۿ<�.�`C
�ubz�ϓl�B��Iɟ�h��y���'$B�D,�y2�U�\�P;��WB�̩r$c��ʟP�	ޟ�':\�	Q%���ݑo[L�Γ3W�ٚw�Cw��'��A�'S@�����?qň�?��O(i��ή�`B��-T|���'m�'_剺i�ĪK|���J��*k�IӍ.(�BH�&�Ojl���IHD�I��l��@՟�%�T�;v0�@
���(T����<78��Idy"���$�6ͷ|"����V��Y4�����dj$'E�rbi�2���Q{8���OĨ[F	6�I�Ed��O�Э�� :_�� ��� Vz����I>��i���'y�O�Z˓j���	��z]X�-ۙ��j�*aL)�I��p���`�k��b>1�	}1�$�a�5[� d��n�IՄ��ߴ�?���?��+
�H��I�Y���O =C$Z�Y��e?�����ýp���$!�$R+V�쒟�q|9��џ0�� �*B��[���SF�ښ^hr�'D�%�Ť�<y!K�̟��I�V�;0� �Yf�HR�9 �� 1,O$�Ze�O
��?���?!(O�a���['t�)�NK�lH���ϖ("�Nx�'������?��k�P��'�ҩͲ5٢}�%�|d�i��)�jc�L���'��	���	����'��AȰ����Ĝ@�ޅ�Bf��Y3e6O�uۛ'BiEBf����I�a���I?f�<�u��*wXУd�;�B�'."�'���'N�DA�q���'��d�_�~-���F*�0U�.?M���']T�r�'un�{��y�'gT}�Ore�w�R
G"��)Ă�����)�'�2�'-�I� nT��L|
��:$��8����BL�yԞ�R$��ƥ��'ɚ-�'5Z�@��gމ�G(�6]
���Mψi|Y`���O����O��Ղ�Ol���O��d�˓p�T�A��Qv�����D�rwĘ����?i�' QӀ�SV�����lĨɷi�<��X���f�J���/yX��$�O���O����O����'��I)J̾9i�y�@�2$D2���I#���j`�)��՟� ��.�l���+�]����Ď�M����?���}��e27P���;�6��������#LC>�
pp %͟t8�ɹ`�:���<c�b���	����Ɇw�2Pҧ���o����ԯ�~����D���kyrlK����'�L�����m��+����3��6�n=�����I0���'"�'�2T���хB�����f�n(�U���S(G=�D�)O���w�'��͂����O��D��������-�ȼ)1ˈ*��D)R���O���O��O�~q%�Oڮ�9o�$M�^P��-0�tJ�'�`����?Q�L����)�O��X�����sLT��K�1^�i	���1��ʟ���ß$�'���Jd�9�A�z��x�4gC��le�Ԅ6P��d�O����O�쫇�'*�V�θ�� �jv�N r���H�*>>7�TjR�'��'��ɐ8��<�K|�����GKH�K��QC�ޛW� E��,����bpԸ���D��%+�yG�ȳ2��"�ć��ҙ*�)����O���5M�O����OZ��쟠˓2/���Q�	�h8
�jg�� 
�p�Q��\��?��'��[�c���)+��
��X����WjU�o��
?c�Xl����͟�����Č9v4�@�?B'ꤒ�@�i�"X$+Z�($����0>��1�P����5_��Y���
0�H8�b�i���'�ҌV [�j�$��)�	�Ĳ�H;���B�g�^v��Y�.�)+�X�?�.�U��?����?y��� ���3e��E�^4���J;�?)�Zn���#\��ȁ�O��L�l��S {��AK"Q8)�����^7��'�Tm:��ѪL��P� �Z�v���X�x b!�[�^���;Ԥ�;duBW�A$U�q:����LR|�D�/
n���O���"  �DIN�0g�ʮ6�N�:ҁ�#�?Y�>rL!`��?�,O����O����O��p3� �0HI��ή"w��1F��O�d�Oхh��)����T�O:�'�F�:0��7Jl$�@��Ԅڔ�'	�>m�"��	�n����D�ˏ"�� ZUl\�<�;`��M��,Q�$E�u�/��O��I�ȓ=�p�T�R�	K0����4}Ez��KO� Ҁ
A�,��`���u���QD�C�Ϧ�Ȗ*��L���)���t�1�߃z�zpx�O��%���X`nA�*��	,�9��Y�a.�3�>����$z��If�Xv����,ۘ���"�vR�����B){�����8V�dȱd��I���Z���
��Y&�VH�!H�b8���rn][d���F�8#K4���O�����5��Ш�l����O�"����Mb�R+<R�z@��/@���3����6��Ƌ��m��tE���� a?�$�ĂfN*H�vJ��'պ����?��	L�3ƴ�Z�ǋ'[`�q:�m��|�ēL2Ua�b�#t8�"Eo�%�	�HO��be�O`xr���5�^�AեJ�2���X�F�1N�QG�|���IΟ��C�Z��	؟��㦅�eO],
���
�[u�u���T�#6���Í�r t��&�'8��s�%Ǩ
X�觟�I)�j1ׯٱ#p���v϶E+#oF��=�J�L�6�g}�D��K�X�J�-�����fj�> �����O��~�'��'�i�&�ΥʓJ��F��'f.�1�Î[�}�Ҥʡ7�Q�/O���Ux�Ex�'�y�i���#`(V+�!��{�`1r��O2l+�0ܮ�d�O�$�O�ҧ�ؾb����w�Ɯ�G#	7\�u� !�"�NP�ܴ[�� Y��=4��*��'� ��!(@�Jr������.�q�4<_졑�O�(f J�c�'oD�'�D�� Ð셺 �.80�4�:��ӟlD{ґx�H��f�Ht%�0���x���8��>��T����\�V�P��łߚ{�SAH�|�'��|��'��	�A��M��%L���QFjE�����\�U���:�ӛ�?	���?Ae���%���3���?���:?��*q��R']B��12	�+r�څ#�g۰=a��Z3G�@{�-C����BSIV��P�Aя��y>M�e`Q3�ay��ߍ�?���|��&ҫ}
��U� �v�����?�/O�$%�)R�4Cf��'��r��x�ra�X��4D{O5�'+�>�q��Bu��K`*�',������pg�6��<��IǦe�g�'L�^>�2��V��BLZ��H!_A��@)�-Nz[��矔���$��"��,2��ҧ�EB\�5V�%N
4�:���$!,1�B�<��'��b��5�ܹE��Jޢ=�L�J��I��zAт$����'Q�����?����?�M|
b��Q��5;�i�c~���ӂ %�Od��<��I	� a��ЎqCnD����Ɵ�@��T?���,6�$Z5UҔ��ٻ�6��u'�T(�Ae��	k��IԟH�i>�	�������ϟo��T ]��$KS�����ʳ#����@=��B��#h��elP�Ǜx�Y��heÐX��$Q#�B��cF�MaZ���N bW(�[g�''"}�'�N�p"��"E��i�!r�ܐ���O���"?��~2������8z��8FǶa6�
�
���ȓI�p4b",ʏ
jZ�����i��'��I T�r"<�G��<Yݴ�$٠�\�A��$`m��}����p�'B�X+�̗�Z�MK��?���i�6�+���!�s���E�<T_����+w�hP���'��ػD��q
�����-��9(ݴZ����ɍisR��۰=�J�0�%R�ݨ&ů�?y��?)����?˓�<�1"�)u�蠡����T�����D�m�
H鰡�_]`�0�V�w�r"<�����?�*O��JЏV�!�6��5Nt�hؒi�B�޵�C��?�����ΟP�	�V���!#���h�'a�%�t�Z�?���eِ�V�E&m���g�Ȩ�a{����ē%⼵"�*�+x��͊�p�4��ɕY,���>�4�N%&�pT�pΟ+I�hY�@�<AR���Z�.��W=ʎ�J�Ǉx�'��Fɤk|���k�8� ��S*:N�jX�yB��#u�h�Rs�'��_>���� ��%��a���:u� F9v)br��	W1��	��@Xf��>z���3}����׌Z�ҘZ6`��`G��sBa�1��'�B�9���To��]�����.��h�ц�5��'�l����ȟ�K�(;s�!�$��w$`Y��"O��Vϋ(x�P\b�Ñl!x��'/0"=�Ohf�H>����d�[��H��E��׆CF交@��B���'��O�:Sp�'���'��ʈ�~r�������x�\��wQ;��iQb�Z0��I�\E����7C��p�%��:7�����M��|a���j�.O*52pY��j��Y�xCgƏ!>y|ÃJ�@㎑�Di�?!��ifZ7M�O$U��Y��ڄI�,x��T��F͙}�p�����.�?q��c*���YA(�tɳaN�<���O��r5f�"��|�'&1�O�B�v���� �,�@��k@�. ����7z�QȒ'�Od�D�O �D�(Ais���O�@�]f.ŸL�f[��G'�;W�����\�+�TZ��'�z�a&CXμ����A�M�2��2�J�r�
G�@��4�����u7K��HO���N
�&((Wi����aP!+~��	�rW�-�޴�?	,O<�� �B>,b��񡅆�ik����̇�
�}Rh�<IF���E/�pȕN��@cHؾ1DF7�%��>Y*���<�!��4=�* �ܴ.�҉�#N��p����){���'�b�'�(H�@�J:��<���R�*'v��1�i[v͒%����`�N�T/���
ۓ6�~ ���ah0oڍZ6<`"\�F�-�s	�*kܚ�����A��{���0鑠2���tG� g��O���<������Z�"�4-��|Y�؀ƃ��(���G{e4�'s8��Џ��<Q�T:E�V�v(��37M���y�]�t�!ְ(���ޟ`�O�n�Z���t@,ɷ%̠W����
��Ñ�';"�Qv�,ys��'��D�Ɂ�~�ո�镖.-��Ѧ��$D��e�¦$��3H�B$�ZK���P��I�m�*|0S��-rSn1���[n�O�<{��'ϴ7-�٦��IB�ӌUn��:�@�B7�T� X�[J��������	4x���4cA� d �r��Zm���V���	�7{��'<��W�I=QuR��H5�dZ�#�Xټ�;P��ON���O󉝤x����O,��x��h�u�<��1�ƫJgT좂?����)#}!ɛMU:#>��"A3I� %��f�k�ҵ�2� hO���>�$�>�%�#L��u����a�ّ���x���'ab�'�\E��O
 en�C�K��%8C�%�c��l��InN��!�=zZ�J�c�@ʓ"9��(���	��n�
��y`����bu�&
�2dBC�	�k6I �MY`RJ�(v���B�I�-v
}�&��OB|�H5χ#zT�蠒GT��T8�.R��
�h���UfTxXS"$D���r$��?��T�#b\)@1���&D��J LW'\qTPS�f
VI�')D��0�H���}y.T�-,>i!S�$D�0�UFܟg�J8$*��� 9���!D�pi@�E�yrL0�2U4:�8c>D�\��ٞ9(��&�Imر�Pc1D�0CɊ�x.��{��^�r:�}��.D������e	�1�����"%��D&D�����[2J�{���,0A(!� C*D���� �4׌�!���!.ʔ1��<9V��~��(��a���{�J�SiM.R���4"Oʹ�/ը[�A�F~FHy��azB�V�|8�ĩ�Ep6��G��Ƹ'@��$![���VO&j�Y�Ƅ��uy!��y8u�MČEh��C�?k�����?�0$�C� e�0rr��/4��!��%����$U-u�2s���b�^B�	�����J�;d#nѡj�w�z���]2�1O��� (A.] ��7��7�\c�iC���x� ͹q,V�R"\%ZfC]+A���d$�ɲ)�j�sCJƧ{4�dG�I��C�I+f[�<A�O��t*8��c(�82�����$��"~�"V�<	d��S�ڎ_C4HI�#�:�yr�T$�����5Nw蚳g2��߻j�a|ҥر����1�2:f�J�MҒ�yR�֑>p��"�"3,��R�f�$�y
� �]���?j�J��DT�bP��+��'$L�J�y��[��ۄ�L/WR������y�ɕ��maRH�X�~�	��T��'>ی�T?ϓ-d���#(1\8�v��6p0�ȓu�"\"d�G�4c8uK �R��lS����T��%:{\]�)�b�`-K�*�?Ow���>�����dB@�!��1c4�^$_k媆�?��]3F2�˓��S�Y�d�H�G�`@���Z/B�'N6ғ�'j� �Oz��F�V�칢 �
^�A�c�G|�IX؞�;!��&���"��U���2�@lӦ7�)�P��'&k�25��t"�l�?����nb_�|b*>}��#A3؉igŮJ��E�&P4�p<i7�I�s��["�,i������,��<�Rm>��U�jK=Xf\����H�I��O���"�i`Q�X�{�Ӄyx�� &X3��;F� �Ms �O"b��O�bĻG�� ��}n�&��ٚ��0R@l�q���w�*c����	�[�65r���8j%Ru�rhC5m�:˓��$��l�2���#6������\�
 1g-ʢv�
5��+��q%� �$9g͙>M�lEcD�ݡx�B�ɕ/�3)���n�D�����O`0롲�6��Q5���Q�j w�0�̎���!�D	5,O�i�o9�I<3�$hbm֤I���*���/T�.�+C��%�hQ�THʬ@ܮ��=!4E6�� 
1���HL���w���1O��NŌA�ș�^� PJ2e��/�8�$,��
m ��9���1B +&�ХK��0�I���<��6QL�J
M�R�g��l�a��s�ޱ�4. fw$�Ă�RF�7Z?-�O�i�BcL=!z�఍�����s�'�(��A��1m@
� ʊ�x��<�F��_�4�ք���� �LM�����"�8% }bE��.�ĩ5��|�
��- �>���Z*޸ BQ%	lB����F�`�����.����� �;C�1.�,�d�z��'��2�D�(8�ѻZ"t�"��dW �z�8b�����6h.7j=Z�ֈ4�PU8������,;Vx�j�*E<�a�B=��Ҧ�A��
cc�!'(�;�n�,k� ,���5=>%��B�?���!��w5"q�����,@s�-B�P]��'8����$E�H�2늅3-�b�N�5��� )^(��%��W�9�O<�7�D�_[4��O~c��
sn~��@�,������'�}��4j����� ��`�F��SCX}&֘n���Apo�k�6�a��T#dd���	7��(����<�f�4ʉ��b#<!��.h��1Rϕ{9�ъ�(U�f4���a_�0p��.��w��h��.�+��q+#�$���� )�hª`�����,J�A���1D�,��Q&�z�T�B���%L|�;n�F`�q.�Y�E�Ә
F���!������� X�)ˠ[�u"�(�,�p�
����B������������ 84Y��]�y�,9k��W*��qëL�@�*��d�]m~,z�a�>D����f�	�7����햍T\�4Q%�nR�H3-P�m�d�`��T����x��X��ND)x�jtyWZ�@<� Oȵ�O���`]	Q����Ҏ��3���PD��iЅ0%�
�m�U�O�g�.�:G�ʱǢ�	S��P�'�B�*���gyb�;?md��S�Ki��(��P0Z!��Ӄ�Ƭ<��a��K�#�U�ߺ>n`��K~�]�5ր��c�,��g	�Lы�N�<<���~y���T}�� p4�����`�Eޅ/����O� FP �ѹi������<�� O�^(��CTJi�����(�U���O�%��A��\�^�kr"O�1q�M�af�RRM�!BB�	Ȣ�i��irLRJ�A4�>U@�"�Л&���1��:�����m<Zk��kр2�$���'d�M�'�Zu�vc�F�|%Y��:^�d�T4j;���V�:���%�I�^�I�D�r9�=9g���>��9�N�$ �F�$͟o�'*��I�0��HP�ğO���z /$S�Y2ł�3;ȱ�ܝ*���Qb�'U `TQs������>-����ψ;PX�x��fp���i[Z1�Q^�\��f��X]$ܳ�@�y���3E:d��%��?,�t�ۢ�Š34��(��c�ށyv"OڬCL�JB�lAqɋ0!�ڼx��M�2��T��K�� �̈g=԰9#���u�%��3�m	d;�7��R�\�v���22l�4]�a}rD��i������z� k`֚=r�J8^�	�!���Ph�-X1#ª�����r�p����'d������B !	n���F	�q �,zR"\(Y5X�R��^�ؖM�4�5P&`E�k*0��iڶ������ ��m�\�	g��-�F��.]�`�>���M��]�����@�hE�$���I$yi�,���I�-cp`���}b@�<�&E:�r&���&�N�f�;{f�Eyԃ
!e�h�`ڴa���pGo�:+�pD�O����z��8����!9^hA��OR�"��b�D��o2��H!;[bU���O���� ����
M��k�J  J��И��ۦm���Ȟx.Z�'�ax�[�X���l@i8=�gHZ��ē��hB�/52��7�E�����&B�U+�O4�a1!��p�I"���N�@`����x�b��q �܂w�$>9V��,K
!9'b�my�K3+)��`@�?�͓gQF��;`��k�nE)e���$#A"�2U�����1��s�D\��f˜mE�tY%�^2X����
mBd�O�1��E���ԟ�$E�|��H���{@`�"�p5ay���.{�����*N�h��	�>� ����s��ȫ#�ą0�(d�1�@+O<���D�
~)N����M5MY�%`�+e��'��� �� S�L���������	Z֞�����/^L���j
"8���9�Oj��B�/Ib� ��/~e����W�y-�7������L�Zvc>���/,?Q4�E"{f���J���w�gH<i�(�?<uĹi7�_�BM�l�Tc�-(:��#�tA�5#�DMK2Ū��3��m�L�����5������aQDq��5����EE�æ����+Sʎ�3�)�l:֢�=EMhe8 �I81�r�ڠ0���:��F�E�d��'1�I'Dw����'�l�P��0}�>x��o�4S�2�80)�-W�}F-pD$Q���xB�M�C���k ��\���ED,K��Ƀ	"�j`��. �Ӻs��D��bǲ�����j�KJ<��<�[��'�b��NDJ@5ї�P��FUp�
6?y��Y�z+�������}�j,gQ�J_�%���S����?y.O�8��Ob�?���j�.b��|��c����5 U��ejJ�H�^�9V�p8� ���-.���r��l܈q	�>х�Ӭ�	�?A$E�^��Fō�6l�]�|
�jG�ܺ(hď�*P�8��$Dax���ܴ�y.?����救LҸ�rl?���ΓPlV	�t��'����ӟ~:��t�B�3�R�05��$W�ȉ�4��Ol6ͬ>���[,T}ơ;WL�W���1���#�~".��<�'���9�|�<�P��b5�}#@�H�Id�8q�BC�<)S��q��&\����c�	{�<����'vl���+-��;�Mp�'��5��#�g��tКR�I��J�@�RGO�Al `��s�[ �ިx&�����8ogt����N��$Ž���?�;��4e� FQ��sa�_&p�\�87�8�y 7�����_4L�u������C3�f�jeJ�p<�@� <
��B����8�P#�o��H�q�W�ii�nZ�E�4�׉?^hXS��D�Vb�v���Q⬋nd�t�r�׹V�`�p��4�>O�]�MXj�2�*2��B(c��6ES1'�v�+͑�yR˟�5&,�놋ތC�(�@�^�i���PCb�k���h�/R�$��7�6��(sG�D��)Q��U�
�~����;D������d�b�j���q~�$ݚ�M+�Unp�(Kd����E{2�M�s (!��G3M���H�m��(OĴ!$�?s!*%��gR�M��팚F	��{w��X�����')&�	5�U'8�͓=~Zy��ɊG,�7
�-�p0CO.�4㞌��7OT4 �V9Rn�`��O,�dڜO��j��3o����"R9�u��'�t,��ϟ�.N�b�.�&��'��X!jR��	��F���^v"�`fF��%K(��&<�y���Y-��	L��L�H�K�LA���T0�6A3�nUr�韱Oh�r��L��E��(B>V��i#�"O�yG��1YZ��PGխL�$=C��|Bg��L�az"���jqcˤ?3X�c��O���?q ���Ü ��_4�X�a��$H�i�O&��M���p�$I�BiL�m�I ���L��UE29O�}Γ��dS�[��̫a��+y��I�/N��azR��|�a�:��6�[�����Z;���$�������(�T�q5�ΰQ�Rc�j�
�=!��i?YB��>n�X��W�m�8�:�˕%%2��t֧���Z�0,��O#@V�0��i�L�>���d�O2,�1�P>�dQ��!S�ꐔ*��F?�7�ia|r(��â��n�(|�
v�F1|��p�l�'>3ܴ��)�1mQ�ժĉ �I�񀠡�*�ayB�>a)O�]+eʜ��]	$�՘I�>0Kt^��$�4o�0�ȟ�EbՍ��C�+e^-c�I��O�Gyr=O�8�$���L(� Y�5ٜ�M��2O�O�g�S�?  ȓƆ�B��Y+p)A�4�N��;OJ!ߓ�~�k/��Y��ч@�8!������dMcX�\ّMB�j��+I.��FD,}B2�;�	h��Bߍh�|YK��)?Tb���5��?��'��ȸ X|6��"+J�*��5�'�F�-^�u)d٫�jV2~��@��'��xx���w�:��)6gZP��'�LU*w.��V!s��X��[�'U�t��E�_� ,y�l����(h��3T$�(JZ�%(Џ@��l������& �-�@ d�τ_kp�ȓ?�\���/�3��9!Ì�����ȓG�д���Q���K��J�mu���5�^�v���5�$2��Ȉ���ȓ7���#�H���a�c����E���d�O(L�S��N_(�K�H� r�m��'�~������jԸ�`gM�/�Fp��O֬y��.}�r�O�(�T+�9��
 #�_Ĥ�A�'�
l�Ҡ�<jbh�K	�Q?�` �O��YC �)ҧ"o�9�iܹ64�s�\�X�*�����X�ZEI7��HQ��)�!���p�xG�є��x�σc�p��� d���aUn���y��ςK�$Us$�R���1D݃�y"��7L�=;��DL�p\��
��y��_n�
%h��Cj�y'�έ�y��O"]h4�Gd�� J4ζ�y2E~��٦mV�P���鞋�y��Y�;��N�8:f���e'���y���ڙ�@�V�D/��AP�H4�ybHA:G&�x�R�@�92��j �y���3l`��vC�E�y��Y�y��� 
E����L�3�b�Z�#ҏ�y�Fɘ<�����!
`\2K�y�k\9b�f�ӓGJ�/SƹZ ��y���1ӧ�լH�;��ی�y2eҭ'�r��%a�w@�X@w�J�y"��H�(�!K:ne>Ԡ6G���y"�-�X2d�BdԈ���B\,�y��"%��+q�E�[�x�V�݆�y�ExR}Yqm���UO���y¡.C��@����J����umطh��J$�'���ņ�K��B�I ���x@�'":5���I�l��X��L�r�T-q�'� �wIǉxg\�Yw��/k?Rt��'3vh�E
�������_��u@�'��ݸ5�P�^u)�n�8[����'1^,��!�l�=녌�$N��|��'�
Y�$�������LY:H���*�'J|͈�%0ұv�[�	ip4�	�'PZ��2��.FYY`�� mU��'��(�ˮI1D,�F�%D"
Y��'�z�˲�ݥwX@�E�@F��'�&U��nD2���*���61E�Y��dF��k����9� ��<n��$�ȓ/mv�IAE�ع���S��ȓ4˖��7a�T������4wO|��Mdv�	�b6}&l��-�0e����l��P1i�˒Wl�:�(���(D�8��C0c�&5I��;H�Q@�%D��Y�*�5�Aۡ�A7'�A$H#D����V�(�i��[����+�>D���E*P2!�� ��@X�8���R�`;D�� �'�3w�z�q�X�-����j.D� �rΛ��9�eW7X��̢7 7D�� ��Z��<~U̴��J��Z��0"ON  v�ܟ�|�I�[�5�2�c"ODx�0�'fˢك"���e��m3"O�)F�۵orq(��ڸw�\�`�"O���"ډ�IQ�;�^���'� pc�ǫ�0���Pqj�*��:��HaB�=����F�r[�~2L��^L�W-Ҙk�̵������'fZ�P�EŹ!����j
�*�]a�S���R�"�>-��.�tQã.��>��OM~��YP1}�����+��9�1�Ԟ|�O���	"ztЩ��G�o��p�����'���[�E��u J!Q�@L��Ԅa! ��K�;�tB�*�(������1�F��p�]���I�9���gTM��dc���*[(#>���8z��%gA�j� �դȪ����Ĩ��5�b ͊��,Or��xk6"�5;h�uA'�ڏc���Ae�?[�jX��)I502��:b�'��TQ����x�ܘ�UC'.`� �\5U*�I�<I���v�D�h�)�73.�	\ Y���6M����2��,��BZ�|r�t�
h�ES3ck���T�x�R8��%��16&^�+�P��)��?V��S��B*g��e�*�#sF��)�ЃB����g�_\��o���(O6�{���j���c�(���W�dqW���,j���"JюklV�b a��D���7f}#3�!L���)�BB4q��|Q%h&����S4$:Ц8-wйz6ˇ� �
Y;qIS�C�:��v��'3|	ԡ 扉#;l(IP���Wn� �\1r����g��6B��(T��!áZ�>�V {a3<OY��i��@҂���g�6�b�!�6�O6� p)�7J�&���	U#����O�-I��I˓ˁ�B����a|reH�_�� ��"hZIq�I!m�8�L��, ��6�5`U.�+���t-�9Χv�x�g.1��6Hx�����5C��5zӇY�W�<yQ��x���������$�<�������#[n �ec��<aT�+���a�3������6Fe���6�!�� B�(J�hT�|�BmY���J
� "욂F��'�v?Q�@p��a�$u`H%_�3fݽK�Z�o�KZ )Z��'��ܹ�Ha��lgA@��̘a]j�)f�"D>�e���9@@�'���@w�v�K�
��j=�5sM?͚�\����I\<t�JaZs�R?P�����> n$�Ë(��4"�i�J�ꇃ�z{�Ł΢D�����ŏ:0xM��T\̟�%n��Ec�] �牕8�-���Ƞ\�`�x��F�#>�ϓ�E�������b�	k�����$�`P�V
N�!�Ԉ�(<���l��DXBJ�t�����#����(�%	bE��J��	���U�$���r1�#"�z��,�%i y�e��<$�br��Dij��OII��2��Y�J^|B����0?SF@�Z��FLR�
L����d}ɜ4jr��SlH��j�,Eo��J�*�=���j5�����ܓp�W�^����s)��2���#ZDɪ���2=���2��#�ޝ2�I��n����@{�*]�|&���y�-]-̺|��\ h-*��e���?�Z�
R���7�R�ȸ���x7�<�ӄ	_c��*����A�L�qo׃Z͘��1�I<l��rQ�¢�z�q�۩(l#?!㌔�6���痛�D�f'�6V����G��36,�!���"M�� Չѯ�$x9g�'f\Ң�05bVax�m^3'�Ԙ �'r�!�f��f4p�A�9"��Ѥ� U��`z�eN��)/0(���I+
���34��;2
!��8�� ��	I�4�g��[5*���Ŕ�a�n�Ӓ$Y!=�
)�S�?�{�)Q����'�i�ұ%��͍�*^�%�	�+΂��7�I@k�$��D��4��P?|t,�B�'�C�P�/����A�RN�0�t'��m���yW,P�qb��b#�b��$q5��;�y�.V�r��mc��V08;ޥ��i�����U��R䀷�MJ<�0���]�
Q;���%<����I�<���g�ع�'L��6���=x�P9��̧i��$�捜��.������1��,H��C
� $��7oq81��ԊPd��HS�9{��S���	�m�������i����P�͎j�8�h �O�%Z0b��q��T�4^�l���5j'�1s?ONdK��׆]��Y�r��1�0<��/ӂupA8V�#
k�@IR��|؞�q@i9h��Q�3O�Ev��k� �8y�\�⃣ $r@͛eo�v� ���ɹV2�H��Ȭ"2Lc��m�Nc�D��nˉgY�4+��b3^��4�m��L{��� /8��$��~
H�2��1��Iʧ�~H<	�Ƿg<��G�6~0,څ���`.z}y�L�0��`�c	ӂ�?Ib�Ƶc4��K�V>� �>�b��$��Y68�T�X���T"O�pD�C+��fLK�υ��d���R9oe�,��DZ�ѰI� )�8���� +F��&��i� _���%i���%=��		Ì>\Oک�uA_� ��1�#��<���BE.Ԉq�����X���G �
dB��,Zf`���	b8�� Pi",Wd�h��W�W�?��'/
����P�*�B�회Z����Ӫ�'#�N#��jf�� ꔀ�ˉ�I�4�[��ެ�Px
� �رD
ջ"�.	k� �.u{"1JϜ=$P�)&࢟���'n�x`�L3E��Id�$��w���1�Ή�9�N!�T�J��#�
I�!�?3<�1�UfX28��8٤�� /�-���'�剾� �����0v��ޒp�6�롛>�`��b�L�����l��Aլ�~�'M��d��8"L���R��C)O��R�n4%y|!��Ŗ4f���їZum6AQ���{�lHa��'����2�D]�]6F95�.��O�/n�C�-�!ㄑQ7�B*1xџ�z��4��!��|��"۬�|C�	� �p"��Y~g$�ࢃ[�t|ذ��A�'���@��..��}�	�ȕn
lpC޷wp���&�O����Z�n&�Z���(��G�0Һa 5�U�֘'Z�@b��E�r����B�x�'�&3�ɡ#���u�4T�q1V��4!n�(G\�'�B�:p�J�<�B��nF*��/O�b�FչG�pՐ5D��>Ȏ���@�T�ypG-�M���:L��?Q'%�8>^�l���Y�	eK٦E��w}�휱6��S#��&�Qa�&ۚ(�Z���fD���I1�W؞���-C�?aA��uY�`��cM04^T$��CV���Z�?�~��%�MU0�85�;fT>)Xo���%��h6H[��E{2�	����O�@��On���[�1g�)�v��>_��QV<O��wN�O���wm�=%En���O�@9 �N�oC�I�/S��1BO�hf
�K��e�N6mZ�x����\!5�8����ũ2߉'bBQ8�]�T��~޺p
 �wU�ygϚ?UKM/�8��'����͆U�*5y'��/M,C͆�P��mZA�"�ć�T�����b���WB �����uĖ*ch�tq��"�O����Q�J�$0V�0�:s�^<z�t�BoN1��!#��D ,�`Bq��r���뢍μp�󤌀[����!�2U���9G*� '<��8�UNЍ\^�B�
1�!d�>�G*תB�VHw�Go��pR
�<i�d��07~�󒃞(g%P��C"�J�'ܥÄ���(:�c�#IK����M�<����f��8���8��'���0\��±),Aݼ}U*\f/Raq#��	\����+�O�j��M1=���Dd�,j��2��Y����)l#�[�K�R���J��i�����9a}��3�$a�s���2$*3�MI7$���� �te�=q��
EmQ���<�pE0#My?yҁ�8��$�ٚl��� ��U�'מu�3FT� �z�.A�4I��'��SË;?� �!l�	]����f��u0������XB��ұb�:�0<��G<T�	�s�ɩKQ ����ԟ��GM�|�����((:H��O$}r�|2`ʂ\��s`$�=?%*�96�б#��-�	�'�~�P��_��
��"��,g$(��%�G,e���OH��$�	)
�|�#2�4�2�,a�>\�bU&&`��$�RǈܕD�4qɶ�_�	t�Y�E�
��������M��-�>�&ыc�1<�*�0��Q���� F`��6����.���B��	�EVB0�(��K�Z�{�(��@z���	�]��"�3D��'@�bW�U�L��%I?<��I���
[�>�xi!f�l��ȷ��I�`�na[Ӈ�>X��e��fj̘ ���u������3xdA*B��&rHA�a���2�O��Ĉj&�$��+�|�;"��I"Gc	���92(ߘmf^y�ē )����xU��˗�$ʅ@�IArr�ۤ��jvz�P��T�P�4P�'F� ^�┨I�P��ӆI����䄈	��R��æ	n��d�����c��3���h�iN����	 Ύ�u�ۭ��"�U\� �g����'ѮY�P�98^�Î*:���O>�˞
zj��劕O����MAyr�O��(��T�\���`��~ȐM���ت2�L�8�-2�m�)<O��*���l�p5����)JE�Ԭ�b�����G#[���.O�b�d�T�Φ��Q�=�ޙj6�r��'�ݐx��2���8Q��>9Z���/�~�F�iܓ_��
�'{�iC82?�������:�ԁґ�K<�E�d?~>b�����X�aQ��Mkj0h��Q�����آb�qO���rdA�%�YQ�I��u쀌��xBiO)���jѲ�<������HOt%����F{��A�`I( ���V�D�V�*a��q�Q98�=��'Q)%���"�;ga�����
��x��v��1l� vF���H:,9c#�PC`h�
m�բ��ɭ_���M�+��(r���jh���i)�T�R�z(,���a�D�@%��L�mU�ч�	�L@$��|�9�L�/K�Fy�L�5&n�CGc&�O֙�!�Y�� QȑV4DY�f-ܕr�#B%�OxE�`!�C��i���,r�Z�)᚟h{Pg@	e��E��9j~���,ʓ ��iyToP)%i�D��*���'ل�:'�� ����L�	5Tb�E��3@i
ģ�l@��RG-��0<��S�,���ۆ��("}�$ߍh;0dɆ�ؚ-����&j���܊��$�{'�tqE�ʂ5�������2#r\�sOJ�"#��51偉�Vb�%
���2�����'f�Z�s� �Ǽ�  �3��L)'4�*uI�E��A��'���P��{_~���,�
��q8��_%6`�X��{�;p�,����'Y�QJ��Ӊ�ē!R�\���[4h�X!ڳKB�j��G}"�ݵ[�D����};$e+��	��?�r�ґ|��e�d��<bP�{ZGʹ]�p,ϙ;Y"X�4ǒ8Tt�=���5c��Ei�KD�U��@���#v���I����ȑ�}�i��i����PB�Jf�K��8��.Հy�&p�OX�@��G�x���*�3) �Dȃ�+БyЁX?�ܕ)�H��H���Iڦ@:�B,;�j��¯L`vB��4gtư{��[�sI�"����s�L�	���D;�,@[X�;���4'��#>G���n$��W�>~�)��Cf��`��#.���R��r����(��j�2���N�? (����n\1*�٩��'��
4	�&zߨu�(�%�����{Ă����B�E�	�4��B���?�O��!�K.=�:��M�Z�PM��'b|��$��90$�䑆f�-Hj
 )$�2��G�Z>)�ـ����H���	=f����¢B����p T$G#�C䉌TbY���
�r����V�b��B��2ʹɰ���{vx)J����"O��q��!"�ڡ��<y�x�"OF�(�c_S����!X�S`���v"O����r��T�r�sd�d"Oz+ ���,�Ar��
5���F"O�y9�L<I����FU7ES�)*`"O�qc���x����$R# 7�m�"O~�A��N�?�b��j�1\<JT�"O�}��ć�j�.�"��	xCa�6"Op�$B��#��B�,�+-=���"OH�15� �t��rm��)&�}cC"Ojm3�2%A�!X��N#s�r���"O,Q���@~:j�i�Lԯ7�ʐ0�"Oj��vJ^�@�h�(F�Ί&�t���"O�!q'�>�r���F��e�$���"O.�⤨K5vhq;1ĕ4j�9��"O�DѠ�ҧU�ĭ��C�w1v��"O����ƚ5|��h�̍��Hj�"O�\���E'H��#Y"��{Gʇ��yr!ڠh)iX�g�U�Ǣ=h��ȓYx��3I�4}���U��T(���ȓ
ed�$IH�)�
�
�&&Jt���Nlv@�v�X�d�2Б�#�
A��D��c/l���ɂTu��1�l�	�dȄ��VI���4!�pq�,�lj<�ȓy�r��¸${�PC�"*���T��Yѐ�Z^T��eN@�[C��ȓ
�&��/�[+�m���U�Y�ȓ�p1�uBNW�^`��l�$���z=�/�2�%�����VZ�(��D�P�%��� ����2����ȓx��iIҪ<x*���u@h@�ȓO��k�A�V�ʆ���Qm�H�ȓy��A
a�ٸq50�b�+@Ԓ��ȓv ���آY�b�!`�����8���� '���D7k�4t��vl�xqGB�Nx(��Vg-*���ȓ�$X���q>9rB�b2��ȓ,�f�e��Q~����P�c9Nd�ȓT,^�������Ce�!��ȓCL��aH�@�0���%v���ȓ������N��DIס�0x�ȓ`T� Q��T`N����A�o,y��!;I��ބQ�,��ckZ����ȓZ�&ICюY#��}�6�O� ��ȓ{�Z����J$Hh=(����p���ȓ8���*�άP���L�c�݅�@��$(�+)(����U��/��Ѕ�S�? "��D)�
B�E
�,�INY["O ]�� XN&P��B��
x�X]��"O��B�F�t�4�B�X����"O��	G(R�#L��G��* ��"O�`��ֵZ̶�Q�	?KĤ8�"O�Z���j�F���QG԰�"O��qVb܇a��I�u+�1Q8�Q"OT��+D!�p�֤쨸Zb"O�	��Gb7xT��,5�]�"OB�3�ռux�!q*�p�@"Ot�iԅ�{�Xy0C�P7l$���"O�`T$�J�p�`G�T�|�b"O���e��E���-R�w@�"O�D;�H�XB����w�8��E"OF�C�a�4���˷;��y�"ONl��n.CM>I����h�1�"OXda�B�>��(����er�e�"Ov���� �eP��ԡ����| �"Ol��p*X_w�H�@TP���"Oҭ�1CL��49+vO�{�$h�"OZ͑�⍺v
Ҥ����;!<	��"O�Q4N?/��sr�))(��"O"��eV6&����GM�3"�bAS"O�R��,7��'̗�X��Y��"Oh���&)�ܨs�Fi�n�1�"Oʑ��kY�A`���
F<,`S�"OlHKS���w|Z�	�+'"��X�"O|�8 ˃�2C��j�?=��Q)�"O�1��Ժg��Z�D�~8��"O^��׈^�/p���ȗ� ٤��"O���B����������X�|Ҳ"O��1�N�f2ɀ�.֮oހݹ6"O�tu%�#/4a���ĭ��"Or]��	D%���{T�Mغ(i�"O����Ez�0�j�-r�l��"Or�`��y���!
ޯ8��q3p"O^�ȶ%S5N��ui��F���"OF<b�ڕ�H���ΐ�s��+v"O����%P0Q��AP'G���y��Iw�O���G��^̴A	s��?>9ޠ@�'\�=��.�N�\�"���~;�Y��'�y�G���QgaV*����'�,�b6���-��5�6�ԫ�z���'��B�0=8=� ���m��']4��u`ʡ
ךeش(���'4~M��- �!�5�䊙�t���'�N�y�&�����C�*sD� ��'��	�2b�6� qR@L$u�Y��'}p@k�'�(*~�|� Ã�p�v1��'Z���I1�2��F$�3pi��8�'�=c�H�HʘhU ڿi�ޠ 
�'��V�mԠI�IX5iAv�
�'XL�#j�Fq-��	�%e�s	�'�쩓g��3*6��Э�)r
�(
�''�J�,P�^���g�vB ;	�'�4����Iz}8$P�fPވ��'�8A$�7fD\R�f H�L� 	�'BR���FNq��N��C2P��'GV�+1 \�b�(m '���L?�D��'e���&dI�c;�ɋ��8vb���'ͬ��k��kFV}c& /�����'z|�:�bٞW�Fi���?3v
��'Ք �fn�(��B2"�-�x��
�'2ބ�`eK�G"Ɲ�LQ��(Hq
��� LZ��?���C�iM�Y� 
R"O���K��3��ҁ�Y�U����"O���t%�/eվb��׺'�Z��"O�<��CL�2�� ��fX)��	�"O(�$� /Ҭ�T���f�r��!"Oj���Hšr��و��:`q��G"O⬁�
�m�2M�5�B�t6���'"O*m�g�S?5�F��HQd�\`�"O�|9��K�ܼ�%'�r���r"O
	�'�,���)A%Ee�dI D"O$���˧����0/�L��"O"�U'�6

�H�"������"O�i{rJ�3m�hq��A��@��"OT�f�V~�@���-W�>)�b"O|��T�oO��)W�;��	��"O�D�`i^�/�:� a#��i��[�"On�q���M�:�"�{�2(�"O,�!��PFj&Q�ӈ�"=k6"Ol��'�h�r�+��9d�Xq�u"O��qoɯ3$�V�
1Ʋ��"O��QCHL�R��l��.¬Q����"ON�w��O�>Ƞ@n�)F�rL9�"OH��h\?w���q�>@�.��5"O��ru�!D���x�,�/w��Yb"O��c���^ڢ�"���}�X�)"O,%2�B�\��L�M��5Np��"Ob c�!�P�
��"�:�Pq�"OR$Ѱ/�qH"��E�/*^�(�C"O�Q7�DB�,Y'g2��"OHp�ɞ������ɨF�2�*�"O�,��Ί b$���U��(P"O6e)#�HdYȜ2S�A�k��p&"OT<8h$t�@�E+�67�\$yU"O��i�D�.<$i�Y�Gg��&"O��BV)T�:�|٢��D�w[��Y�"O J��(i�������9@l �a"O����c4ߪ�:��K�K�i�"OB��d*�EY\yI&�	�R0h�"O���b�]�d?^�B�du�nH��"O�	�b	�R.>(۔E̴i�@8J�"O�x�*�NN�Y��
[?Q�"O�
����t��X1uʼ�V"Oԭ1��ưpv����@Bp�ļ�c"O���n�=��n��@��0�"O�E�uJ� Z�:���"U�
�"O4���#�> �-ܥF0���"O�H�D0PH�G�X0�c"O�4#��%��@c��SK0$�"O�Q�4CøG��%kC܃1���"O���E�8�1��ᙎ)��m�"OĹ ���!)^0a��BD�S�"O�	Bb��
�A"0�T�K���b"O0w-3ZjP�j�	��-����"OL����Ǭns�� �֍!5� y�"Ov��I<'���Kb���� M+�"O�p
���%D�x��ަa�f��"O��å��St>V�i�qҩՙ�y�
S�me�l�d�\,\���6�y���G���P�M����rJ܎�yrζa6�aC�osR:u�5��=�y�&GAp�}1e�Fq*�QrЈ�.�y�)ؐJnC�=1��ī�)�y�l�.'�0EЕ+0��Z�hͷ�y�j@�1t�9��5�ʝ��y
� |=��� 'X��T�LF���R"On jg*g��(�EO�Z��5�"D��I"�G"=vиڢL�	9���W">D�H�6+��b�J��ŋ
k��U�D:D��1ի��]��'JO�J5s�#&D�(���/�2�)7�ƝN]J� P�!D���R�.i���H�{��!D��Qf�H�6#�(��ɄO@(��3D��!�^�ӊ�isG�=hrB�"��2D��b���j�H�_-+Ne# /D��xqLҔe 8�S��[ ;���@�*Of�����0<"ܐR%��tg�9�"O�L���Ħj/����yc���"O"d��㚴m��T[2i�*_���"O
��U��$�A���85D|%�&"O*պ�h�NXzeA:ސXK�!D����";�<�C�%/cNȲ�?D�8K� Ь_�����{4B2��=D����a��;%��� kFO�.(P�(!D���1P�"NP�@5Ťm�Z�P��,D����)�X��X���69CNA�O*D�@��ƽBn�"IN�8�csa&D���A�9���*
�o�X�Õn?D����A�p�s�>�P	�O=D����c��b͔�0A!��@��-�<D�X�ӡ�@���JA�x�ve��5D�����
:���q�kӾ5BF!Pn2D�A�C[�a(�3B�;_��lJ�k2D�ԊfaVR&p�a�J�*�$�k1D��Y�`��~�B 1pg�p���XB�1D�(�m3Y���$���y���/D���&K hH|�h�Ar�)��i/D�� ʈ3��0U	A1]�`gK-D�d�&d_?����UȍB&!D�٠D޷r���c��D\]�d4D�4�`�����]��/�7�N�9�2D��P��'z~�Ʉ/Ŏ$��#g+D�`h`��1�X#�E�.����'k)D��bq'	e9h`K�Ą>�<A��(D�(���b�ވ�#�X�C�xu8�j2D��k�*T�*"9Y6M��R�F-{si,D�\�գ�*���pHY�:)�F.D�<����r�Ѩ�K��R x�,D�<A %R�-���q'�	�v��tM D��B�N�s�Z���<0�N�a�-1D���Q��+� �Qk�!\u,�a�3D�� [*fB2���c�R?6���5D�,`�J�Sm�ع6&���t9�a�3D��9�ޛS�Az��̴dFL��`n3D�HK��͒�.H7X-vQ���>�!� �}<b�ۂ��B�%��G���PyRNSX���h$.h$�3���y.[�)%j����0]p���喯�y����r�n��4@�M�y҄K�~�lD�����(S"�]��y"dZ�_��ph��@��)'�G��y�DA�K̂�{�%��C�~y�fH���y�& ��a�)T�;  ������y"!�=i6�8�#��6�Z���Җ�y���7��};���4/澑)W��4�y�%���i����<�Ԍ�$B��y�D� a�uF"�/b`jc�K��yB��(b��`z4Y�a��)�J���y핍,x[ׁK��L�����y
� Vq��Mφc�~��Z,7(�`�"O�م�ÃG^��eO\dh�pi�"O]�����T�L,�A�ޅ_���u"O����N<`q�@>��Ș`"OXlքۥ8�u�� �vLn�ҧ"O���ኵ`(�1	#�܍	��qY�"O��,J1<r��Y�DQ�Nu4@"Ov%�f㉸K�ȡ�E�vb(qR"O��B��tȒu҇E��dXx���"O]�e� �>%��ꎷ4:��k�"O¹:w)Sni��"�ڑ��i��"O���G ���/V9Tp�5"O���+e��DE�҉'����"Oz4b�Ŵf�n�(�.��vٴ�c1"O�TH����2�E@����"O�i���P�^<�0`�N5*�CW"O�M�ʿW�й�����"O� �ŀ�4�t���ː-v�p���"O�y� �9Nc�$��J��_	�=�P"O�c�ʙ�,�24ct�S�DMh� �"Ov��j���1)ܫpF���"O6dCdE�v��#��I�M�$E�"Ov���"�~�xb�%�4n,��2"O��@(��-���wĘ�oX��"O�a��'PGE[A�5b��q1�"O0�!FN�.,)��*r	Q'��Qa�"O�=����r���r�v_��Bp"Oq"���x吕��͝Z-���"O�� FC�u�dS��Z�H�@�"O�\�q�זfl��5K��In��cG"Ov �`{�X�L�WS���"O@uB$
N�Kx�"
�
SFNІ"O�P4Dի!�@��!ɂwV�����iH<a��"� �IJ�Q���5� _����?1��I%Z�C2,�aJ yJ���b�'Eay�OZ��&��T*P�(E���CR*�yr��, "���G], 2$sg̑��y��Z:Y�\�JER� }��-�Ν��Bpt{�̘7�:X�4f�:|H8�ȓp������+>��(ץ�<$�h�������F��&1|aH�d��3�h���sUv�s�6y�
t�`���E}R��ue܌����/q}�e��)�8�$�Dz2�'k�(���Q�|p����<Jv4�'!�%�q؈LPz]+Ъ8��s�',��ÆDͱ>v����Z_�|�	�'�R-�C�͎h������2��D��'�"���2!}�	q��?ʘ��'��y�3"�Q�TL� ���:\�j	�'�-��`N
 �N��%��-1̼�0�'$��g��]g��0TM	%�0��'̾ �뙮C$�Cϕ�� �s�'���S���ͺ1������'x���q�Z�EŐ9����dR�'?Rt� ���Vr[$c�$�.�:�'��9���q��I���$��0��'��{�V� 3�뵋P׈5Q�'1� u�#I�Xٰ��:3"�Œ�'������)%����k�1���'��q B�ۊUbH�Q�0ܥ �'h�9�e(�#^-r��p�
<�FѨ�'s��pȑ#�H���D25$L��'�&9ʳIE��dI�l�w�����'.�a	�L�W/�4b �
o��4�ד�ا� �8�d�fCtYs��'�4�K "O2�q4f� ���)��G��yJb"OZt��%XDr���k{&x!3"O��%���l��yhr)�;�4("��$1LO���� ՛5!�c��נD�~�R&"O��X5aP�tQ�FՁ��a9�"O�	1Rˁ#�����Hl���'��O�!cU%���� S*a��"OĽ�2���c�����U�tm�$��"OFt�uo�+!
��%��4[ln���"O��0����B8yRgF:vj�}H�"O	`Ђ�K�pR���7�"O�ɧ���]��2@��-�:X(E"O���dh�F�¡̘�`�,�[���7\O�u�h	����
Z�@�q�"O�㢋�9s#0���+]84D���"O �1F��C,j�ە	[�g��"O 87��`hW��y��a�"O(���_^�}�2���k�b��$"O�I�/�:u�@(��D��?�B�3�"O&$ g�ص9x��y�L�8��Dӧ*Od�P��F�x0�%N�ln`ъG�)$��� }�غ�(�0A�XP��;D���"ϟ5h� �1c���&���#e6D�����%f�ԙ��N6t �o?D���J��mFTiڌ��B�'�C�I'q'Z�ڒe����eI�
��C�I=%ۀ��Fn�? ��`8qjߖ:�XC�I �Av�R($�����a
�B��:u�����͉HĚaО��C�	�3j6M�b&-�,-���1[.C�I����q�F�]��؈�c^�4u�B�4r�p��ԷK�L��c�<P%����4�ɠ}�A��D# ���U"�~x>C䉷b>عp�źDP��2w�ڌg��'�ў�?u#&�`3�Lc�D�5!ᘥђ�<D����,��'���uC$iZ�	!!8D�Dz�ː:|�v�^,sp����4D���K�6�B��`��g�B��Em1D����8:$Ib�(��G,T�T��]���@ ���2p�U`�"O��H�OC�|̀ծP�sB��p"O�T1@-֕5����犢T!�#�"O�ɢGk³%(���׍G�R�e"O�����Q�?�hԩr�� d���)"O��C�����)��QZ����S"O��e��!
�pH�qEӢ�D=�v"O8�1Ə�}W��� ���Knf�S
�'���̣nY�KQ��./լɪ�'�J �5O f�zͣa$պ#���'�� ʀK�]������R(�4y�'��3����$QI&a�W���!
�'�|sCA�0:`��*��T�N�Tmz	�'>"}ZĞ�[�vق�.�/Aq6� 	�'�Jii�Đ�H���;ū�b^:aI�'��M��L�[�Դa���U��
ϓ�OPu�t �ZZ�|8�S�8�ڶ"OF)+3b�>&L�@�J;�4��xB�/�S�'TQF�S�l_*{��c�As��L�ȓo�<��©^�v�h1����u���ȓ&d�͑W�I��2�B�����`)f��9��LcK�?;GX���D���O�6b�z�H�oF�x@ȓ8¶Y�b"��$�0���ƈ�/Z�H��S�? ���6e2�Li�Pꅬ|����'"O����ؒBIޕC��L�,��"OZ�!S�I��"҄P�&����"Op�s3,L2K?Z�RVb!:���X�"O��.;!��9w!�3ȠE"O$�v;S(!����.T�@"O,)��O1uFl���E�?(=D�s�"O$|K�jC�+f����#i8��"O����V"�M�_B��R"O4����� )����LV�+��Xq"O��q��6K⸡ ��V<�0�"O|m�t�\m�d ��¶S4:у�"O�Ku�� ;7TQ�p@��c "O�1C����i��IZ�J�<P�l[�"O�,���X�k�t81R�r�d�SW"OXh����1Eڊ9	����=n��s"O\PQ�KI�|,x(b��Ì9RT�a"O��y�-20��p��Lld���"O���ci����6+K�b٘�"O����UxxP`w�ג&�����"O8�ɱ	��)XЍ�UI�s'���"O��U%�>�������p4"O:h;1M�>f�\1�o���"O����*'�����_^>��"O�EBt F�[z�����#��Ę"O� gJX��2X2�Ȇ�-�4�[!"O�L n�(��9�8j��
��y��ŏ`I^���tְ1��L��yBνA�2��,����u����yҦ�i��(��l�!I�L;����yˏ�!ޠXhP���u�Õ�y��7J����%�T��:����y¢�G$�ܨ�������	�yL�̲x��� ��FLV�yr
�?N��8p��rp��C6�y�Y�2��jU�ۦX6�Ycᓝ�yRc��:|(�A�L�L�P���y�n{X���(�<�+@�U+�y��ɬh�"�:$[2v�<�'�M��y��QHl��s�@�1����ʸ�y2d�9�.\ѷM��*Zx����y��W0(p\�s�"P8t�쬢!�ԭ�yrdǽ�:x��1g鞉`1�V��y�!_.*��i"�H�t!RD��cٌ�yN\7y�ض��
u��4Q�����y2�@ E��X�wM��m�e2#���y���>Zf��@,wʰ��ù�y"EM+>��	���o��Qa!V��y��MC���T�@Vk ��yB�5��9��K�%j�`�BL�y"N���2��'��![�l��y�O�N�!���ɲ����֜�y"��	ڠ�FN�x�����y�
�$V��lSD�_�&�4�q�
��y2�2�x�bE�N�;D�K�y��q��,�cč+Q��`���y���/Y�u(��ս���k����y�� �m�`P���T�EQfp�%���yB��
L�����7e� [��I��yn�/*�܁;	4x��y�����y�ဘn��e�sa�B�H�)�#�yr��"Z[���pe�@��,�D���y���[�D�٣a�
8v������y�!��F����b�9��������y
�  ���X�>��Q��	�r�N�`"Op� ��I�$^�D��cB�E`ʀi!"O���?pn.����$sPɒ�"Oz�;�%���6�O%ghٳ�"O(L0�C�:��_�I���"O�y��ņ(��k��û[O�i�"O&a���.>`YPՍ7��p�"O�	�i\�~n�����Oo�h:�"O°��O��l�kG�mR,� A"O�Tг�ާ
��D0� ��OH�!B�"O�TJģ�z; ����-*�"O����픪u\v�!�+�,�Бp@"ORa�qW�K���ˍ2_Tp��R"O �X�� �GA�\��	�06G��A�"O��+kĵZnl�*�N��=0%"O�`��AJ9J��)d�C�}5@S"O�4�c��%$�s�N�I�	"O.U����/?^�A�T�@P9W"O�b�/T6�i �EX�<��P��"Op�Q�\� ��IIP�[P�(�C"O�EE9�ʘ ăY9-��Ƞ"Ofmv��m��T�B6��-p"O
ia�#\��� �P�Ih|�f"O�<)��'Z���3��#����"O���e�Y}�qr�%�,�q�C"O�	��>oL�K��͎&Qfس�"O��a���}pT��$�}�� b�"O��B��E�L�jH))��,��"O���әBEz��oX�c�v<�"O�\s��
N@.ئ��T~���G"O��%L�Y�lI�5F��Eg��B�"O���p�V�4]kc�(K��	E"O�i"ҪRm����V#o:@�"O�	Akˤq
��匧'R(hjU"O��� ��©�5G����Q	
=-!�dZ)d8@�噍N�ب�ը!#!��B5T#��!£��A���]�kl!򄄮Y��|�D��$����H�M�!���K9E���=�����h�R�!�d�jD�� lR��m�D@�!_!�Z�hZP�g�~�Kă�XG!�D��d�_�B��!ra��+!��]*�K�)O<;6\p�"R�!���\��)%��:hP�$��~�!���%x`B.����:#�!��/u[MȤ�͝#��p���&<�!�ʦJ���#�"W60�2�b���5�!�dW$B��ed����Ź�L�.!����=���n�%�įV�!򄎍5xzL�3%�m�`ac���{!�D���L��8��A�a�_#Ra!��/�|�cq-6o�u��G�t�!�D��A�0ȇ�U�5[�+s���<�!���Da^L� F�zQX�("�!�ĔD9ƐA�k<ں�1��I�/!�Ѷw)p��æ ]��9��J"!�W�3��$c�|r���K5B�!�D=)i��Gk�~�����7:!���J�z�@��F��l[�?�!�$�.:��Z�)og���"A�5�!�dE32S�y����5Oih���K�!�+	ma���mR:41éF�g�!���[�Z]�%¬|`��Yd��+$�!�ɞ4X
�@gȭ@R*����X�!�� n�����p	�Vf�?x�mh"OJ���.J�3l  �
�7$�,�"O
�HAe �$��7
ĕ\  @�"O�۰�2f� 
D��F��"O0h��G 1��S�����`B"O!a�F@Q�,
=wr���"O0@�t)�4}� #1ʞ�h�Z�Zq"O�	V��k� H�iZ�	y�5�'"O|�=�i�qGߖul�H�"Of\�7B
�3���1&O�bs��R#"O��g��.���HGF��`���"Of��f��XBθP��K|1��(R"O4Yg��Ni�B�%J�Ԁ��"O `��J?x<�C��^�>$K "O��C4�E~�0p`W� D���"O�9C��#x*$Ո'/Ҷ WzEC�"O�US�o!.V�	�	j=����"O���gʰGF��$��V��C"O�l���Dd��-y#P�1'"OЁ��(��Zfi��C�B8E�"OR�x7��J��y��ʊ�|k؈ѣ"O*M �i��ΐh7�J-�:!x`"ODYa'��in�8��F�tU��ae"OPp#�V�v�Pٳ�ٺ1H8Q��"O� �a��`6���&
�99Ќ��"O��t�A32Q!$+�4/8��"O�5� �V�J���z@�]�q#�<�3"O��Zs%��U����8B�$�"O�W�8Fqȹc��N_L9� ��Z�<�ei{���2�產�.!�p�a�<y����8�Ե���R��}�2�e�<��Λ8�u#UL�I��k5�Kc�<��$�J��� W���r��J	]�<�N�`;�x���H $�P�nS\�<Y�fڮ.5���u�$���L�V�<1��\?���D���Z��I��O�<!���M*l�A�� �j~��K�<�g͌7{�P�*Bg�xjI�<�l-��4��֕-"�`�`y�<Y*R�-e��Y4�<Mڈ�C���q�<�D�ɤX���pׂK6�6J��U�<Yu.*�d��S�-�X�!,�|�<��F���X���b���#�+�v�<�A횕#	�����s�, �&
�t�<�����hA8Ԋ�<NH�cp�<� �5j����☹s����%�G�<	V�.u6hm�6�ֱ5�b�����y�<�2�+Ĳt[�ȍ��I���Gt�<�����L�@��C ��D�A"O�S���)�F��V�ɚ9�� ��"O��r���#����e�$f�ĝ�"O���1��7upJ+?���5"OxA�$�\��@��f�}�`+w"O���#��\�qY�{�4��F"O��A�
؟�ҹ�cO�׸9�"Oz��f_0�=���ء~�x�"OX�*�I�Q����G/���"O�I9��F�YI�����2v��C�"O|���x�� �@�hv�"O���� ����"�#ܨL��}�b"O��iG��b|��!U���|NP�"OT�b'�6.�މ�R�6:��p�"O�u�f��c~��h�E��}a�"O���Ѝ;�}���z�+�"O� ��� ��<#�5���a�����"OZ�sL�!v�<l����:	�mX�"O �B�9or�2Ae1	,]�"OF�0W�.%D���Q��i�P"Oh�*��D7�%ctΫ�<��@"O���Oѥyg�р������ "O\�aFo��$��5j�Ȟ/�I��"O�p�Y�H2 ]���9n^y�"O�a���7M(��� W�M��"O�`�\>w�μ�d��?��1{�"O���C�KPlX��Bw(��""OX�Z�<�P,�=��x���_�<9��^^���B�^�nAAf�P�<ac��0�-���E4�\�(XA�<�K9S���{���]`eH�G�<a�̄N�0�Rb���L��� ~�<�w�RY2��IG`�ks\��SCy�<�tJ�$"E
T��J?6�yq��w�<1rjȮe��tA�g�Q}*8	"ƍ[�<ёD�/ .�YBf͂ ���Br�<�f�A��,��`��F��-�ALm�<iD�G7+l��݄b������C�<�FR,z�X�zW뚵A���b�T<9��)O����7K�2d��� �H��ȓn��m���A�oڤEb�L�f��a�ȓeI`���"���t$j�jK�Kh�ȓ[Y@�� �+w�xm���3t��͓�hO?���-E�C�`�g�ǩQ�U֠'D������_��BC"F�ڭ�2�)D�l���RiV��ǩ�6h3�ͪC�2D�4i�I�!��1��:$pQ-D�0�"!  h|zU$��#khe�#*D���',��vg`xa%�Y 6q:G!<D�X���Wg/6	s��'p����cTqyb�|��9O~ذ`��)����u��iO���"O�H� ر���^�G����U"O ���JK���ďx�����"O�z��w��<�����^^�!���2�T�wE��@��q�{��'a�$Y�!B+�92w���|�@�	�'�^ع��Y!T稝���E%o<Z-ѝ'ў"~����te��` � �a�#��B�<b%��Eƈ1����K��� bD{�<����|@C�Y��J���FBu�<A�
�6O�Yi��ܾ[�C*p�<�G�L#�z�2C�M�(��@ӬLe�<��*I;M;<8
�n]�2C���f'�w�$��4�%�ݣbMƧ�zԓъ8?	���n��j��j,�8���	M-RC�I53�nQ��WJI�字��B�I�G���cǈ��N�z+1`T�ԼB䉌&�JѢ)[I6���<��B�ɍ)d8dQ��Q�ioS�h��>��B��,�x�t+�$ �3��*����$�OT�O��FaR�d>�j#���^k���"OƉ�2�5g�fuQ��6pt��a"O��13�I�8���b�3Ab�P"O��1���tB~��F�(wZ�su"OU8&��wY6��b�:kD�a��"O�[�(P'(	F�H���SB�}jc"Oz��!IE�i���a��/X0U!"O�aE���1���Ud�&9����O<����s�l9@ۧS��a9�I$A�!��/P�hMq������i$*ʜ_x!�� ��u`U�P��=k�(��.�� "OL��.U�m�X4ФAX>.�R��"O���Q�jX����7b7��1�"O^$z�ˉ>Xk�Ѹ&��8.UJ�ٔO4����h����� k�l��%_�b��-�S�O�fBm�q�uk��B,�Y��'-$�dX�YG�R7��%�����'7 u�soJ�@1��w�n���'�j�a�fۯy�(�0rb
'����'<J��`)I�`� tرN��}{*�q�'���X�"�?/k��A����r*���'*����!���X[`ƍ
{Ѐ(��OX��ʁ&��e��o��Luhr"O,�Bg�߹sGx�R�ڪ�N��R"O���s�I	0�Hhl�>k�,�c�*|Ox`�SE�.�BPprd� 5�*M���'dў{�a�Y� qH�c�8)�E#��(D�0W͖
"�
�3&�ξi!#%(D���6�Xu�ء��$&��E-j�h����gx(@*���%�\�#�X-Q�pB�I!�d%A���\���Z���VB�ɉ�0�7���6��Q ?T76B�I�*��D;$�L���ɤ�U�`gB�I�F�:�JҦҋi�x%I �G�&|�C�	-��e��`��KO^�q�E�\�vB����qC��#z�,��%cıh��B䉖uy�P`�o�4�&	�t#$y�HB��+z�Ε���[�L!��/��N�ZB�I#ô�#�?��US�^B(B�I>^�0 ���JΔ���^�c B�	&���qD�ԃ<�v��ȟ�G< B��`O<��3� Rv8��J	;ݡ�d��MhY����X.�])RfӯN!�ҊM��C��(HK�S% � zY!�Μ$ �I��äW1��;`��]<!��J�gL��3၄}��
�K��h5!�$<?�`Ur�,-\ �"��C!�D��~�4CIȠ!#�,Na!�����RD�D������?Vx!�D̒�&q�d�ۦ$g�d��
�'�\�B�ǧ>]�@�$Ӂ_��'�z�:�i���Q�D�RN%Fe�'�j$�ƁbW�	ҢN �KU����'���b#_t�Y����Hh<J�y��'��O1�jq۔΅�a�f쨗朼7����e"Ol���o�r�>�ҷ��Tk"��g"O*!	j֞RS�@	Q��p8dY���D{��I&b��[���v���$Ú�I�!�D��	���E�ո@�HQ�S.7�!�䔦K�05��g ,��t�0K�	
z!�� 
T�KE�N���0X�Űuu!�B$5�@D�q��4H�ThC��W!�D�<�(�`�ʣu�v�s�&0*!�Ęk��H[���'}��=��d�!�$��I6���f
U�`��f� ��!�d�34z��&��$$��	� �ۑ}�!��*�ph�E!9e�F%C�.�#I�!��w�(�{�@4yDTj��u-!�d�U��`b��)
c�dY$Oq!���40*J��aI�"{=�HѕMMU!�&�i���Һ*6�"�k�8�!�D�@ \��_&Ox�J���~�!��,x��	�Ip�޸�f�D	kg!�dOB~��j`�6�j�S��!,A!��O� `qj��{
@����]�*� ��'�ў�{����ޫ{ԊB��=g�$)�ȓD# I�b�(c��5t�6|��HJ"���[�i�9�gG��K"N���5� `u/�T�f��C$Ij����8� !�"-�D|�%�
v3`!�ȓdMڵ��0g$��)�Xn���ȓors��[��Z���)&,��<�+O��=�'}���P�܀L�Tt���\!F�"��ȓ٪���`�#:���u��*����02��u�\"&b� :%LR�?Ƞ5��OR�����x�J �� Jm�ȓ:9�Mx��F�h���)�'�?� L�ȓ5d�q3&89�v���(�>~�潄�"��	 5,W�s���[d%�U$vY��?1�B�	����CѱS��]�#)�B�I�	MfLPDB�;'�В�Cŝ<+�C�	'Hp��I�dL䘹��߭H�C�	�p��b��U9q�A���ݪ�`C�I	H��`������t@c�9`DC䉇5�T��cNӗ-[���#
�p� C��ɟxs@BЭB�Z�X�]D�=c@}���IN�S�O<�E�s�Ӡ'�p�H��1t�68�	�'�l�IC�r%��4��y���	�'������nS�����	Dx�<��'N��y����44�u��`�:O戸�'`$Jf�W'<pR�8�c�`��'.�]�fP)2��
r���h��')�̓ee�7?Q���Æ�TD��'c�X L�>�������,�ԩ��'cR�s�FQ�/Z�#yZ���'�3��V�}��Qi۶���'�����@�*�	QoO�
��E�'X�2��P7L dPX��X�}�>�J�'%��A�@<��9�i�x�M��I��c�,H|�Q�f��ND@Uϓ�?a����=�/{J,�
e'%$&�����n�<Y%�ܡ\�{�.F��$�B��k�<)0c�
Z��DKc�n
��H��d̓��=	�d�=&���jR�����f�<�"hR�A�^�a�E�E�T�P� e�<�Ύ���X�f��9W ��4%�a�<�f��)i��#�ů �j|���<A/OR����Y�~0	V�Y���IQ��v6!�dF˶���Ά���@����!��ǡSSpd(�S�����{1O$�D:<O�t"��]�1y�P�+�[崐�"O��A��]�l�"��A����g"O0H��iB�)/�����@'��-�#"O��j���P�d5R�0�6��C��Ie��p����KڀLq�uH�i�E����-���y��-Wm���B�,�6@�Â���y���*���� ;�$x�۫�O��$��<�*˪A%La%�3u�!�䚱j��h h6d��ZAh^�E]!�� O$��[��V�-Bx2���'N���8~�^X� �><�F	k�O�O��=�'!�a���Z4Z<BBA��k��t�ȓ���F����M/|D����'�2���"9T�'HŞ\�2��4 [�pnzC䉓E�r	�6��P��B�Z!yVC�	{	��Ŏ҃B���Ƀ%D�\C�I:a� A����:}��"B�B�	0|v��#�, �t�+M�M*Lc���I^�S�g�? �X*�g���� ���_�`U�$8U"O.��A��J>����L8���C?O�ʓ��S�OZ4m#WH\�*�^�ҰWiU�(��'���a�dM�7K`���H[	�ji�
�'�X�8�
4NR��G	 TJ���'_H�� �.!Z���Y9����'�(HYtIV)�L�l��^��1�'[|�R���0f~9)0	�BA��y��u��`P���~U��wV��y2�'F��|�����cjI&��_�a��2�!�$�1�8�* ������P�I�!� �Zޜ�hQ�R�8d� JqAJ
G*!�d4cj�6#G!E��RƓ"!�D�\�I8F��*?��Ҵ
ӡ6!�dT�l��\���÷�|閉�@�!�@'�b��ͭ��uY�'��q�!���|���.J�R�W)6z!�dX[:�ụ�HI���+�h	D;!�DȵF��P[ե3�&�(�HF�$8!�$�7TDl�D΀=e�����m�:�!�$�]��x,�"�"4�1M���!���-�&�9CF�=I�Fqy��#z!�d�#E�~;�g�d�	�@	�=�!�$#Y8`z��RY����dbE�a�!�D� (��K��6g�H���/�P�!���d�c����n���0%ϝ�X�!�V9UgV����� ���q�!򤉵iPؙ� ��HN�X�LYt�!�d3�"9A��J@\$���[��!���N/E�* C�	��9��r�'(F3'!�x����������'�9aV�N�"�,Y��#_#z��,B�'���I^�,����<�
)��'�qkf/�h��qZB��=3�b}�
�'3��P�kiuƤ�F$�x���'�
��e�ͭX�>����@ʈx�'�!R�A��Z�CՎ$dV�	�'��`��#Ձ�f	�P!Y�>�%��'&.܊ׁH�Q]l\�@Q�}���S�<�2��\����6A��^8��*�O�<i��]^(�&�?z�@�pXH�<�D�38gt�BG@8g�fM۠��{�<�6���r�,� h�B( T$C�<Y@�J6*���Z�C@1[k�h8WDt��$���1� �`I2�B��V�_�� K6D�艦c�դm �� n�$b5D�k$/�?!tX]�uC�/b6����>D�$[jH�U�X�w��L�)��<D��[U��5C'�5"V�T�s��{�N<D��Q �':Ǌ�֏R�r.�գti9D��ISF�9�Yv��CI����1D���4�Ķ��%B#�ݣx����1D���	U���	���R �"��-D� �B�U�K4�`0�����`���7D��P������җ]lAK�9D�����[)�����(�F�APi8D�<S��Ь7�����͚�y�|t���5D��p�âB�B�y��(X�2��4�(�OZ�Oxe�'�%yl����ے;&["O���E���?"�����_6p�G"O�D�n��&�V af�+H��y��"OD��k��N!`�U���Y�"O�D8� �>4Ԁ2S�L�!��rg"O�d{h�.Ȑ��G���)�n��"O� ����=��L�6��Q�>4��'��	�+#��I�@�>�p�r�M�m?�C�I��䁛FRJ�!�V,hR�B�I�'��@h�,��P7"Y+s�;qt�C��-+A�@�0�/d_\L#�Fޱ��C�ɬb��2pP<lV`���ުC�I�h:8�q&G�%��cX%��C䉩'��m6LzD�qv�{B�I�{e�+  "\�e{g��5��C�I;/B��Р�`%��Pv*3 0B�:�H�" K/,b1�W�l��C�	*��4č=]J��"q�ەr��C�I����h�;e]�m�mںs�tC䉳V�<(J�B;g�z���$��6C�8]h��jǋ^D~Z-ru)�7�C�I+`1�(KB��0�@��A,̼c��C��73l� (؅^�E;Å	�L̨C�	�*��E1��[�i�&)����$%�C�ɋt����C�֍ �
i�FR�B��4A(��qB�Xc�8�M�_`�C�I�{�ƍ��a�/H� �§�m��B���"jSSw�\Z���V��B�#H�R<;�Ȟ�Ev$;�lQ"H�B�,*;��9#��o^b�$аk)~B�����B�Qu8��hL +u�C��:&l��$��8j�rI�f�unhC��:F������؁B�=hF�.G�<C�I9�d�n�!	p��)�A,� C��<6t�ۡ!��a�BA�S��6m�c��D{��$��C*8�çϟ�x{��;�y�V5еru��s���`���y2�#?��*�ŔxW�)���.�yR�8[X�(�an��l'	���O��=�O�����B��QZ�H�-��l4����'rL�*�50�.t���J�l�$��'*
i�q'� 0E�M��ϋ�j/����OT��O��O>)s�S�|�P�K�ET�s`�<D� �����W����+��_��(�9D����)W�6n�݀�e-7����6D��4�V�0�te�Oϳ5���VH4D��1��ڿG��BG�M�!M�[)-D�苀��zJ�(��!�Ȓ#,D��BA��`��"�6־ij1)D�0�!��"Q�:H��ѓ�y�aBC�4�;P��@N�;uH
�y�d�)�0���N/,l��D�K �yRJU�e��9R���D(�@I�y���?^Q���6$H9r���"��	�yr�ȫp�6�S��'c��Ak��ybEB�	� �ӉK#��!Y�'M��y��Q�d�D���C! m2p%��y�`I�9�8x� �	�
�@?#�xL�ȓWL���%a�F9>���]8�ฅ�A1I�% A5���7u�n��@e�A�	xf�ZSC�%�ZUΓ�hO?�{EG�l�����*%'�u��A2���Lt ��Ћ�d��b��`����"O�HG���iA�K�UN��BE"OjxT��!tZ�Fj��[���"ON�ڃ��Q�"]��c[�~��mc�"O:a*$aXE���q��٨uv�tk"O8�{������BEѧi�ل"O��7���H�R)����>P�,��6Op���˳����B�S�ʨI�m�z !�� �5:ԥ�=�ΰ# �Ȼ��}�"ORD[�/ܶ'��m�6K��"��Xi#"O �aG׏@�$��*��h��E�t"O�
�oܠrdB��ϓ��@�BU"O��@^{� �3ofHb"Oظ3E��2ZX����pO�Xh�"O 9Z� ΂FP�9H!�R�lfj�z�"O��X񆝷P��kD��|6�@R"O�T�Bn�7Q���@r�]�vdڦ"O��r�'K/Y&~�ѓ��� ��8�"OD���@��X�^�r@���|��`��S������W�8�1횩7�v$Y�Jܓ\�!�ċ�v�(�1*
d��=ʂ*��9�!�d���J5kΙ��Z� ,Y&�!�$���G"�O�\\��[�C!�DS>˄�E��3H�����ӎ"�!�dS'S�^��0��7����U$�]�!��q�4Y 1/E�;��� C��~�!�$@-F5�Aqʙ��jMk��SK!��;k�"��JP�l��f�-P!�Dʰ1�TY��	�}�V��V�.A!�Ā*G�DM�e��(|�Q9%��8@�!�I�`���S�q��9#bBW��!�L�?��l@� ����Z��
r�!�D-4o���DJ�4����a,�!�$ݲQ*��һ}���F!�,1!�DìcZ�c̞�~� �p��ɶ@�!��,q�q�fS�j�H���% �6�!�D̴P+p�Q-E�ܡ�b	�9�!���	td�$�4a
�X�"Wy!�bւ����N[O>��a�(I�!�O�y�Le#1��-EB�͘��Rm�!�d���mQ'��@�;��8"O�R�HL�
�4��TOӃ&��k2"O� ��n��	�8��ԍ�esd"ON���ޫlt�}�5M E��k�"O.%X#C�f�����Y������"O�����L�H+���n�s�F���"O��������� '3�����"OT�s�8>��j�m�ٔh� "OH��GɄ�]��x�QJ�)�d�W"Ox|���l��ǚ
@�E��"Or�WH�i=R���D�@��"O�d[5��,��=y�F��#<����"OXi(3nы=��u�e^�7V�1"O�����*"�dH�'1�L�a"OV�
eؠ�3v�ɜpֱS@"O�I��OK�qp*u`�mޠ:
�D��"O��ip.��O�YqW�	d$��R1"O��3�D��A+�%�j��x"O��$�����Zt���_���5"O�{�b�<.�^,P����X�H�V"O����]1u�n#S�ӫr�%b"O�B0MkJ��T�1�y�T"O�Ԃ���X��ź� �;F� "�"O��)�\�^��d+�O��6��H��"O��$A�!}�4p�,T�~{��KT"O.�cB�&� \�3+�(^k�,#"O��b�5&@��H���jU�"O�)+�D�o>Q eZ	f���6O��D�����(2�X
�ZQ0���aG!�H	O����N�I�������9^!�͉n5�Ԡ,W�Pa򇌈�Py���:0A.$Bu��E����y
� �0�VԖ$��i�w�G���"O��;�I ?�$p�FߊM@�䒷"OL�!#��\ăd�

N�*���"OĈ�1@��8V�<1Xy�0���gF�<A�G�1��mB���m�P���RE�<�C�C��Ѳ�/ȍ5��\1o	V�<����6Dz����A�v��w��P�<) I�]�T���� �Πs�iM�<ᐠ
?"�Ї�|�wo�m�<т��NP�%K6�2x���CB�FD�<9�A��P���-(֢�c�#Sj�<�$IKetd����(]9<���]�<QjN�
�v��&N�0�X� ࣑[�<��+ck�� ��7~�<�U�P�<���81oNm;q$B�rJ�X���UN�<�̆�_c���B O$N:�K �^�<	���:s�����;G�H���hK`�<a����#��Q��*6gi����_�<13�ӬlƼ�Q#��Ѥ�!��r�<1W(ܪm<r)��`MBĨf�An�<����6E��ʂ$��:�R��6̒g�<�昱v&NV(�2�酳X6BB�ɦ[۠�#�u�.�x�!A*�:B䉀-�J�*W�
>Ĵx6���\L�C�T�
�#�&�4=ۜԚ�B��S,HC�%8񠍐���e�%8�a()�VC�	i�������1��3���NC�	8_��2�M�/�#G.C�39U�ғn�OL"Jī-t��B�	kQ���r&Au�<�Rh�t�(C� ]�����)Y���Q�"��C�	6E ��1�܊np��w���b��C䉽Wnt�Yl[�=�Bݨ!��)�B�Ih7�4�f�HlJ�)%��+/B�I \���Є$� �j�C�ob�C䉧E���EC�)f5 ����'#�C�I��d�pGkԔ=o��X3L��Q��C��M�>�CQ@�'kDL�ʒ7��B�	2k�Xc@,�{�xl!�nVB�Ic�f	bo�A!�a򕅋�E�\B�	;j�l7��8ot�c��HB�Ia���!��S]N)�7���B�	��(Rķ9Tt#5IŮ��B�	�E�0���F�L5�`D�C#uՀB䉅Ո�:��Y'YY�4��"E#B�%7��=���?%�D���D�Tj�C�ɠ% �ij)W�;dt��##קr�C�	��"�z�C�U\Tp�lV{�JB�		6�\�H��_� )*t�g�,$^8B�I .u��{�˓b��1#m�@%2B�	:r��f�LS� �׬P��B�I0����DUR�R=�ǌ��4U�B��>��M0���*(V}�f
�z@LB�ɺI��-Z��C/g>�̫�	��VB�ɑWb��
�`��p��| ����jC�	|�B�H�R*S��S�k+#�&C� ��2�Zvw� �I;� C�I:0�8�ic��a�Q`E(�'#�C�	�3�0U�e& �����J	*- C�ɮ,�a �ץ<G��ag����B�	s�~�1a��Zb���ǊG�IX�B�WRD��!�k5p�2�φ%D�C�I�g<�X���^jqAHB<��B�ɢ���@cA�pz6��P*��h4B�)� � ӆ<w��{�f�V���·"O��[��ӹa{~��Z�+h)��"OqJ��v�ed[�*^Hb�"Oݣ�"W�O��e� ��O�TT@�"O�dy�.�*�PuA�S$-��B"O\��n_�U�����B��u��"O�;��J�j�R��E�$|�T�p�"Ox��"�X�w
��pa9w���"O��`��E�oJ`T���=ta\٤"O������"}�h�χiQ�$"OL�y�A��@� �?yH̍s"O���ì PY�e�[>֨Br"O�(
�?��`j�78����"O��pT鄩:���6Ʉ�-�r�"O�ɳ'C:�
y��H&T�&"O�m(w�ˏ"' �Wǘ*I08�"O��F��`H-ѓ��zd	@"OD@0��5%0�p�1I�M�v�36"Oj1Fe �+�P�0�f�9���S�"O���p��4c>ܢ��P���B&"ON�#�+
Pw��Ƅ�[����"Ov�B��>y|ƕTf��h���t"O�EV�kn�m"fߙ2���"O<��h�C��(�e���d1i�"OJ�eFɦg"��X��տ �	R�"OfyPC���{�hz��Rs�HeXv"Oj)�G��b;��ڗ��2�h`h�"O|��7��t=��H�Y�xA�-��"OdbPA�<t��� d��z6�1J@"O(�j!��i;nT1a�L�p'౓�"O�����S�@���ju�6&:ɫs"OJTc�f٭4�"���iZP�D�+"OZ�A�KB�&,%�+��T��H0�"O��� $�]�|T�A
	`xF�y�"O�,��8sђ���	DB�1"O�IWG�)r�D]�ቝ{�v�t"O��!dIN�a���FO�����!"On0(���\��U�Ϡk	�x��"OB�P�3��i�l׵�&�R�"O么�D@#-X�
@&<����"O����8X�"lS%�%�XX"O��AB!įx�J��k&����q"Oθ��eG�]���#pd K��\a�"O� %e� 3B��dX�oWb���"O���&��[��#�V�5B(ղ�"Ov��RDD1E��T�� ��9���"O��b&oޔ.t�z7B�p��p��"O���a�eNp����6G�xD�"O�MH��-;4*4�6nϮ7f�t2s"O�t��K_*{��e bL^�<�R�"D"O}���:J���[p�6d�
,x�"O�Z��(d���		u��S"O�!/JN� q�ڇ��(�a"Od�# MT�Q|��G��O�84y�"O���#��$U�6,;a/;HQRAX!"O��b6�"T�����/�t���"OLx�Ȏ��꘲�MAi���"O����7`	Z�l���5{�"O���G� y$Ak�P�a�:���"O�3�D�4D~�쉥,�~~���"O�� ծ.uu4��e�D�.eV	�"OB�4��u�=[ǉ�;U�E��"O>}!GD<A�MCU��G�ZP�"O$�6㙮;���֣ի�,4��"O� �U��AT��Ջ�@[�*�\8jG"Oa��C %��(��� �	g<	��"O���4/	�r�<���-X/vR��C"Ov�jŬ��,��	��n\���"O�İ�g��*��U��RH[�U�"O,�ʠg�P���:�Ө}�D���"O���&G	7�t�9�h
�5�n@Q�"O
]X$�	�am =iV�O�9�4H�"O��5'vn؜���2�T�{"O�	ytdZ�R0��!AZ�����"O�ac�bK�#2��HA6|��4"O�P`�`O`��1�G5r �x�"O$R$�#|�����Q�@=�j@"O��@RaL �i0c40P ;�"O�ȡ��1.����a�06� ��"O(�4-
G^��C��f= �"OPPpQ&X��V��s+�+��Qۅ"O>T�O]�Q2��0PӍh���y�"O��ei e��M '�N�=��y�"O,��UÕ`,I���&���$"O��[va6�4��F`ۑ!��	��"OV)�W�)u@[�N47�T�D"O�y��&Hv��@tn[�ꌛ�"O4U[e�G�����4� ��"O>�#�DU�kOn	�����+����"O,�i�%�&%6�z�/�)ew���"O~,c��mB �`��#r]Nٲ�"OB���I-=Ϝx�lP"Z�RQ"O��%���V-E���MmJ��"Oȕ*@���BC�ybSeO94~8�q!"OR��a�]�h��SUCDhf�P�"O\9�P�,R��r�C<:`�K�"O�%�#'��M�&=�$��l6�X[!"O�y�̟sTdѕM��Q(0�84"OŢU�r֘�۶���|��� "O���L�p:p���J�#s�Dx"O�y�TO��q.ʱ+"E�`mJyrW"OZ-Cƅ�`�A{cيb{�y�&"O�D9fχ$Ƅ�3���>rx�b�"O�!�'�E�QQtԈ1^�fY"�a"O�@	#�B����a��t^�I�@"OT���-F$[�����R�4U�T�1"O*� P�Q�BĜd\A#�"O�ls�,�Z�FY���E�vJ���t"O�� $��#��`��D�H5�""O�arR�ߢ|�0D_3A�<D�"O����"��4]�C��Z���t"O�A:S��*^��SŮ1U\��"O�Vف;-&�S���uK�ȹ&
T{�<�db�O�:9�0H��Cb	��G{�<�3����0�b��;PL\T��/Gt�<�6N�?3�:�R�6���g�T�<Yq�
��4����	k�A�6EN�<ӻ4���@S8��4�K�<�2G�I�A#ׇ�sg�|��ɞD�<	��SFcx��S�H.L��%D�<qD&P�� R!,N&#�L��`��~�<)Մ�qwpi��Þ||P�� Rf�<qA�ΖI��4c0���	� �c�<GoV3o����C��x�&��x�<9�@�C�6�`�ő�nT�=)G�p�<�2�"yG2,�A�H�jk,@�F�Vq�<��$ܗL������2S<ؚg�H�<����j����a͓�3m|]"�G�B�<� d�!j?�t�耒�xp�G"OB��ѭ��xǀ%9!-�Fq�{�"O�@��N%o/�SR��8	�H���"OdR��Z�N�B� ����df)�"O���G��8�\���"X�c|�0�1"O읫�D�o֪ �d�C��`;s"O��p$�>^�(� @�F�ά��"O��#R$&\Z���������"Om����"l)�SL��e�ܕ��"O����k¬gڸ��Ƿ'&�l�"Oؤсj�7s2�EP�l�0-����"O4@T,�5���"1�ùg� �@`"O���R�@0��8~l�I�"O���D�^9��)j`oـU��i#"OX�h0�ϫ5��x��Մ�Y�"OxJ��s� s6�"����s"O
�!'��G���d�����Z�"O��*��%z�ctC�@l�a�v"O� �gB)N�2t���]?e\��"O� ��Θ0�N%R�cc߆�sA"O8�Щ�5��B�ዯa�6�S6"O�ip�%P,XJ��p׆�m�6��"O
��'g��0�VP�eG �<�F�0d"O`�{sET�z\�eA�x�FU�E"O�iV�[�B��`q瀐��:�"OF���*����%��b�c4"O`�C���9d�\�c��,���"O���	R$|���f�3,��y��"Ol-�U�I��L�,�	��H�D"OL�s3N�8n�Xe�4��v�JM�"O�Y{`Gȝ~��#/�95�V���"OrT�(�>��p��K�1�r-R�"ON��5�V�H�y!@@'#ښ\z�"O�)Q ��r6��K���) �i("O��"Qꄉb䜽�V�$l*�Yrt"O�99e+ܩzB`e�T� (n�h�p"O$9�NK�O�8͐ң�3F�٨"OD�����	�V���F\����"O�S�/�+�q�ğv��XT"O0\��%V��
���3��H2"OB�B�Ç&4�LrBl9}��d��"O~��Sd��p�(˳J#���"O�����߹��� �F��[��h�"OfQ���.h4�K�7���KV"O01��'����$�8�n�� "OD���љ�����#�(r��@!�"O`Dyb�8��8ǣR�}�d`X�"Oz�`�� �/e���v%�/9pZ�b�"O������01��b�nW�%L<H��"O ��C�U�n�:��.N-6��x"Ob���>�Ʊ�𬁧t�����"Ox�2(�a��m
Q̔7�y0�"O�ZtF[�(x��샄?ũ "OکaW��1�H�1+\�\��"G"O( ѵ�P8z��P(t�[ ���b"Op��B�x���2b�s.R���"Oh���!=(e$Q@�
 ��"O�1b����(-�T���(��1�"O�-p��W�s�ā�s��:$��x3P"O0��ʡV*J��%eZ�
�Ĺ+"O��QQKOe�&t��ٙ�R k�"O���FΕ
:1��)� ���ʐ"O��5Ì]�+5'��:�r-�"O��5GN�d8��r��0W"O� *���*�ggzlC�"Ȥ*:�ܣ�"O*�{�G	/:౨���DX�a"Ob<����fiPو��ӳ]y�`ҷ"OPK��R�ir,,[���^� ���"O��관��oC@ѰZ"�0&h�y��Ȃz����釸$�u@����yB*�-ld.�:̎���98 "�y���27Z��"�
a0I͑(�yR"мC��dSb��(�&E4�y�L�	CV���.��3��P��y"I�')��yt��y�4y�OU.�y�M&|��2���$O��Y�����y�׀C����e��Z0�����(�yn�dz�SuB�9
H�����X��y���8��!�1 �N8�_��y�֊k��8�w��qc��a��1�y���
�$���	�+a]�ɛ7m��yBkȗa�\�q�n��_�1:'���yB!��s�&A�4��,W�N$���yB��gz�e*7a>��8V@�!�yR+�G�.���ԸYz�Ȥ�>!�D<$~N�q�
,5�hL�tOΕ4�!� mx+���;�v��n߸2'!��,6�B� _�=����L�L�!�D�(M��;�e]�!c؉���[<�!��	�Tܜs�%ۻ.�N��0�1G!�D>�37!L�!�Dx;T���Y0!��8�	g E�z!y��K�!�DQ(\SJ�0AM�NXY���)3~!��@����p��@�.̡�l�7@!�D�}��YC�Rd�RAt�A�F:!�=O �J *��Vɜ89�jP.:!��;j�\�0�U7m�RL��D�7!���;�X|Ie�!��dɥ��w!�O )�<�����0��QZ!�ݰ{^!�� $�la��*oJu2k��E!�$�)3P^U��Q�[�x�3�(d�b"O$(i3ė��L �Śs���1�'��8}R��@��1{�mV�E/�� G�	1�y��V�4 �) l�S��h�1N��y�6brف��؍ ;����_�y��31�@� #�&O��0=)�"!�AL\ӥ@P@����y�ˉ
Ǿ�1����^@{e�~��'��!�oB4*�*P�¡+dݲ%c����0l��Mˠ�@"PO��{D&�,&D:C�Ɂ@�lBp�=~�VX���Q��B�ɞ=�dI� M9:,��h�]'�B�I�Z�vu�E��3Tq�#�Fb�Z➀D{J~�9sm�M�%���K������b�<����jk~�!1��(}?0BE�b�����剘LM��;�k��q�l(� ��9q�$C�ɑL�F��D�����@K�f�~� |��)Dah<�kK�s�V8{Ac1|P����hX��Gy�)� p2u�*ؘ]bpi�����yc�x�la3����X�r��p��9�y,���^�)��(J�0{q��y�c�q�� �a
�TY��� ʍ�y�#!�Ma��F>OG�<�(��y���1ZN��CUN��q���E.��y���VeR�K(�=l���qv��p>�N<��펏1O.Y����5�N4҄�M�<Q�#NW��KW�ˇj��y�B�YG�<)��U��d�v�
�VÒmFc�Y�<� f�#�^m1��S�j�`��'�ў"~
����~M:��e��?�����,��y"���D��b�X�5a�0:�E���y������\�*���Ƌ2�yre���b ���?K��a��G�y2����!��[�N��k�/�yN�)Ue���oŨw�]᳠/�y�+5RF�" 8eN8��#�.�y�& ������;!fѫ����y҅Z�`�T���G[��@5Y1��yRLYFԡ���ѩ��y�S憲�y��{j=�PJ� C���I��yr���.�[a*e���"����yjP�E���OYbx��M�yi�<%I��@�O�X�P,�3�yR��|�Q���X�o��Ժa���y��Ҳ8K�]: c�=9VhQ����1�(O�����"2xpk0��O<�E#aO?,!�$2��Y8q .a�`����(O��
O�@)���`
�z��B�!��n�t���:X�m�V��$!�g�B�`��#����lģq�!�d�H^t1�@ƕ\ ĳs�C�!�/)�\[FL�x�XM��9;�����w�\M�������[F�+Y�C�I�g� ��d�Z��u�2g]�	!:�ƓFUF$��J.������:����� �����<M�h��BY�xp�ȓo���3a�U�@~*��=_ ��ȓ.��e�z'�� ƣ<G������=+Bϔv7��d_W[إGx��'A�Tb��P$#�r�ɡhҰE&N5��'Z�6*^:L3��!���,*�MS�O���d�q��xɳ
�-8PQ ���a}��>?ѠF�"2ry����$,�e�g�<	`�T v@��s��
x�Li��Pz�'�ў�H���a�ɚ~�x`�S�ڱo�D���%�!q6��3y���;Kí;�T���hO?҉�]:$XC��$�<����<D��F�]:]mP�3Q\t:S5?��+c<�Y��V24m� �&�m�HŇ�u��;�lO�?�
,ʃ��$?ڨ��O ȉSw���kR�Y�!ԄA�Ն�w>���듫<�t��BP�,���	���	���o?(94.^F���p�*U+#�*[i���Ќ��h��)�� 0"�`�cڤ!�=uȔ�e�t��� ��1�E�n�FXQr���OR���X��P�`�%i��Q&�V�||셆ȓ
�%B���ye�ӷf�**��x�ȓ�`���$��q�)1�J}��#o�E��Y �2+C�f(����^��M�`�Y�o��Lre��Z� U��	�~=O�Ș!LE)��A�	D7qt�r!"O����ǌ>��@#\��E[d�&����O�6��Ot�#���w-4�C��^�uB����B1x�d�:�'��E dO�~U̜3"m�x�z��*Or��O(��O.4ꧭ[-h~��C�e]�>ᐰJ��'I���ZX��P�+W�qED�C�I�zj��T"پX�}���;Q��B�I��)̑goDH�1�]�B���:�pG���ZX )P'�4`�B䉹�6%��gd��P�m*E��B��e�@����7Rd�D����z+�B�)� ����L �P�`�kŤPP%r�[d"O�y`���-���W�T0�i�"O�	B �~\��DBD���"Or��5FD�-�9���R*�la&"O�X��	��)�$86!�b�"O�H����"���Sޒp�j	(�"O��0`��: R7c���R���"OD��j�d� 1{qg�r�ޕ)c"O�dҁ�߳_��H�P%�;5�p���"O�1�u	�%v��8���H�:�*�O�$�:<�p�S#�F�f�,�Z��;E��'�a|�k��|��X��E:W��:@�G7�0<���$ƙ]�΁۰�X�s��X�2���Re!��K�P	X��W�D�l��c@��~Pџ�S����L�L��ZSRR$#O@:2!�D�+�l0��8~���#nY.>!��V���[E��FB�1��'U0��xr.�>YM<�ێ}��Y6�]�4nv�9���r�<Y��WN��Ո��Qx0�)��gr�I[����O0ipń�C�jSO� 43�A9 hV�<�4j�<�4��G ��-?B�!fQ��p=I��L;xP!�v
�� dL�<	 ��8@�� B�q�JH�G�E�<1ЁE�(�S�<�,zg�YH�<�憙��X�I_�Dw���A�<1��*5���a�mC��<i1
r�<���:4 jUI�%N�1Ǧ�[���G�<yt' S8��"$k� +3��]�<	7���C�T����@d���a�<A�aտh�`�S �^F �G�e�<��Z=X�$�p�C:C�t�PQ��`�<����Z���z�b9lp��	���[�<A��9T�)*���-]�p� fWn�<	��O�"�µc�)^-)\UX�$Bh�<�@�,y01B%ϯ{�<����e�<����1 �c��I)ʔl8uG`�<�'g�$�(3�C�f�BIHC�Lw�<Q"�$SҐi��IC�_l��$�Ou�<yQ썤.[A�T�D�vHt 8�AMy�<�U靕W�05�䪆�)[hu0�ll�<AgOK38n�-����5p_6p�d�Ni�<���μx ����1S�(ȇI�h�<Q��1T�-a��l7�e�Ç�l�<I��I��Ā�KXܕ��)�f�<Yq�ǁCh8a���?��H)�Ki�<y��O�����iQ�:�<��jQf�<��R�Q�@����;���r��i�<��*�9�^����$^h�Êg�<Y�+U�Q�X��9(]�T�E��{�<gnڧ8/�akN�7P��� ��L�<�5���UX(��W��;	�(dS�mTF�<Q�˙qO�4�S���c@�1�5J�<�� ��8)���;m�4�$c�`�<pe�?k��d�@(¸8��$KP�V�<I���<㈉ ��-J氤�P P�<ɀM:e\%H��ګ1�|�ʲJDK�<C��]�x]�F�ьMnZ�,�E�<ATG$K-"|�	�_����G�X�<1�i�x�Ba��
De(Qz�#O�<�.�5rJ9��ނ]�$\c���a�<Q�F����	�E>.��0��C�<AǁF�@�F�(�`�T�a�T�|�<Ѱl��`�u�G�G8D ��x�<�����hh��� 9�YᡮN_�<� &m�d�]�q�!�$�fBP�[�"O�]c����<:X2�� 	=�(�"OP��f�
p	HT���|}���"O�	�F٩u;~u�7���D�6���"O␛Ѥًx�R �#��$�TY�"OHq:��,�22WA9V�f%��"O铓�I������۩r�6�[t"O:�p�P�@Q�,���G�,���""O6��fš(��L��ɖ+]�e"O&� bJ�DWp]��(J�pr�K�"OJp{�Nݓcb��F%@�����"Op��sK `���/Ȭ$r�"O���F۷Xfd��&������"O�y{��I�j�H�R4�,,3P"O4�jD"I�8:(���?f���8�"Oęz!%ܲ/oa"W&V�zd��c"O�=���01�e1E	1)&�[�"O6��S���2`�‌m�A�r"O�J�}����#Bm
���"O��$���� �E�8���&�_�<I2��Thv���+ "g
�0@s�<��/~���{�#A��
,q ̉t�<�C
�l.�Q��b͠4��rc\s�<����n*���u�T⑀ Əu�<y�d %j;Ҝ�w��9�� ��r�<�wi�3*d	XSn�XQ4{�d�p�<م�C�u8|��̎�:< lK�,To�<9A�̯oH�Хc�`~4�"Ǔf�<��è�f=�r`"33��`C	n�<�b��������J!>W�(�gn�q�<��&[�v�$sF��"DT"�SW,�n�<��Þ�m�r��*�!?�\d���l�<Y����h�ӄ�{���Ie�<9���3]z��R��.���4��c�<qF��_X�%ɄBG6�����X�<��J�QHHq[�͑� �\��-LW�<��ެU��ЇO]<N��͘u�I�<I�.Ѯkט�7�5k hD`/\E�<ywcԄ|����t႕/l4�E��Z�<��Ș�4zLC���2BܫǏ�Y�<)G̑ ����r��iX�����O�<q7�1�J�R �VG��a�J�<�"��%Rﲄ��A�B�A��A�<�'k˘A>�- 5L�7SZz2�Wt�<A"ꆥ[�6���]=^48
s�<��n�
GR؛��Ì/GN̓e��i�<���R��Dʦ(Nf�6,�1*�i�<���d��`Ӓb�0ՠ��N�,&��+$��V	4ݪ���'&�0�b�*D�<k��)�Lbr��h�tr�E)D��[��ũ}���:�J�~�0}��+�OԢ=E��1%��p"��2~�x0�Α=	^!�5%� ���� ��zy@��=G�Ip��(���J&U�5����)�32�L � "O$�Ka��z^m�#I�G&�c�|2�'�JU���#�$��q��L��'@x��0DY]��DH5&ʊn������|�OՠH�n��P!����_�U>b<S�'9� �q�Ԋ_����A�?Vذ�
�'�|�'�I�8����� !�	�'�bЉ�$��:><��O~�>���y�I5lO�<y�&���Šc;���u� 8i��}B�OZ�A�	�.",y@����A��ς��y"g�/ɨ��D�HW�&�ಮ��HOj���H�� έ�g�׈A��q[u
R�sJ�����'�Q�����8QX��w�T�!c�4�4��Oj�=E�Dfv�H�"BM%&�2��"�)���Q��|z�(S�a��)r� s-p�I�� z�<�5E]&�r%��L;,�1�n�z��P�'��Y� �*��0��-=nܰ�'ސBխ�" ��b��_-ʼ�'�"�B$`�ʄ`(�`�2LH �	�'�m�W�-X�����'7�=h	�'~l��ǈ���A���"�����'x��Dy��)�=�&l!eS<K��+e`Y�j!�$*�dɇ�/�pL�@�^�IP?A�{��>1�O���@O5w�f)��@ >�i��'O�Γ �>	P����8�	�M�U��8'�H��ɤ81mBG��E��ʗG�+�|��:ғB�f|��i[�6�2"���B>Vl�'PڅDy����d�<����y��q!ŀ"��)�\�(��iP�hԴ���͛{x��O<�
�d�P�:��1���(/���~؇��r�U��v��(G+c����'��*vo9�M���W �,�'�Xv���W�!YC�ӽC�.���'2�viמYxhL�cC��%/��ۓCА}���d�O�O?��@8B���Pb\�|;�c���1�ab�O����A�f �6��Q[,`�"O �4��>T�<����|X(����p�>���i�.@�4�n�7?x1�mV By!��*Lժt&	�(�.�Ȁgdf��U?I�'L�b>c�ģ��-����$�Гw����+�hO�ӍB4�$��OI��"@�S��6--�H�)_<2��P1 �#1�� �(�O���$�������b�yu���,B��R������߿�D1����M�"���;ړ,NV��u~N�R����U9t�ȓv�D40�	ѽ~�"ɺ%k#H�H�ȓa��j'$����V�Ýv깅�n��8!�F��8��YJR��=�D��	q<�����#sԠ�υ�*z�5y��D��0�<)S��-�H{�i�m��=˒�C�<9��"���$���W����f�؟0D{���(l�F�;�k�$ y�]IFi4j�C䉷V�(WY�D�����<|x�N>ъ���ʜb���2͸�+CŜ�F��{�D�2T�,Ր��v�p�y�D."�!�Ć=[���4
��.ɢB��Ȭa�!�ĭ_�$ĸ�N	�`�49��ᘟ�!�d�<h��=1�@Ȋw�z*!ئ\�!�D19z����C.[E���x!�dގw������U�6.�5�h��"OR���\ �P�CB��+݀�(w"O:XB��Q�c#ެ���e�WH<I�m˓\��BYJ�t��o��Њ&��M/\Dl�9և���qj���`�!�G�(Kf�����V-.4P&�4L��'F.XEy��4��&�j|ÒJ�8im����#��O ���)ֶ$�y`��O�5X�jO.	5!��ܥ!^@���i0Oڬ��K1#!��B	)o��1�f�jX���
�5�!� 5W��m��`�Vl��AǨі0;!�$�*:1�-c��)k�2�;��['R!�	�b�<89��^X�b�KGAO. �!�$	3f0(*wfڸr���2���)W�!� �B�j���1q�pd�@��!�d�2)XE@]�l2M� )"O� P�)�	E�9**M���g��"p"O���MG������2���w�'pўl��h�bo�!ɖ���
�	�ҁ5D�x�!�N�?Ǟ!�k��&F���W�?D�D�SD�?�F�pФ֐S �1�Ј!D�0�����,Ԃ����g",�㔍>D�dQ���l "��6�C�l��X�g�1�I��"<�����K	�u���*0�\�x0��:�"OM�0��#�*TcaΟ�<N��T�m��?�W�>�&�R�+�N�
f-8��͈g�@g�<�FO��!:�A Z�}�|Xgg�y��-?iK<���Ɇ0�����ˀ�a|��86&�&ba�C�	8&Ѕ@�c?'˂dR�mݝE.���a�W���'p���g.�4	��LJb� ���X�j4�OV扬��4��i�9�"i�6d�

C�I
4�1�%T�B�<Q"�ŸTEТ?+O0b>Z��C+�����(.4���L*D�lK���")�NUy��/=�D	�C-�	^�����$�>@�nԴ4���j1J�R�C�	N����!��f���
C��ʀ�ys�#OhD�*j���D4}Ba�$��,�r��(��+�+���y�b��d��]�nN)�FNO�HO�=�OP:��&7��	���`<��
�'�,�c�GÏ��@3��J..�,�Q�'-�|�e��!\���Ao��-��l��'[Ja�g��?Jd� خ/���Ǒ���'��N?�ę֊�
4
M(H��<l�U21#;D��%.U��z�&@�l����EFF��xr@�ӊ]�Ƅ˲r��k��+�yr�}���Hƛp>h�X��Y �yb��*8�z����i`Α�`��yb�a~�H���a!�H���ì�ybEŕn�v}K%h١Q�����`���%�O��2����cHpvO�7�d% ��'���?7�l�T$A7��HPCN$l~$C䉱'vD)��Ѳx�<�C��'X� C�Ɂ 8�(�kϒuwX�@��M��B䉑D������'���V"��w_�B��s��a�˭
G~�@�lQ �B䉽B���2p��P�'���M���#����O`]����e��p�E�E�M2��'��	�?�@��f㕟|V&��Ì��V��h؟�Ca3�P#g�Be�Ry��2D�胷��+z2*��үߦ;QX����0D�V�&x���Nm(l8�P��yR�;I��'0���si�M�<yE
Q6h00�H,��A�B�P�<P��R��Sd�IW�*��4�P�<)�ʞ�(݆ݻRj�E$��HQ�BJ�<�B�^�� ŤP����A�<14'��@*JTȴdȝ5���ːg�s�<�a�?� �ߤ2�h()�Q��y�R�	��r'�U<�t9�h���y�������1�"�6C��yht���gဋ�\��fnݺ�yR#��JJ�d pO�t����甹�yb�� aw���F�s�|�QHݦ�y"��+V��z��E/^"���4E��y���]`F3d�Eq��T.�yb��,�*p��͙7W�z8C4�T+�yr��p�V���FV�UX �9�%
�ybH߬]@���"B�@�}��G��y�S��r��*�ITM��� �y
� b���*�4��෠	��Ј�"O,U�ł�+"g�q����=��yPw"OnMJ"G��a 5�to� ^2��@"O �a4#�[R@D���D��z"O�����Z��賣�8+�\$S"OpQ�L{-�
ìV��U	�"O���'&�n	�1�B�/�N̢�"O��@�
_6r��f��<R����"O|�K�!�$2��,*ߖ!q"O�eH�č 
�P���:��e"O2�9rNΈF�@HB�h	�?��"ON S�Nо�dy
�A0l�$��"O��K N*U���	�f]�SL(8��>���DW�/��yӇ�I/rs�i� �(xP!���]�ڕP�I�th>d)�A�/?!�D�8;v���S���FU`�A���Fq!��)Da �iÝ_� 8�R-Ȓ2�!�<M�̴��(J�՜ݩ���$5�!�$�[�
Ѡb�\�V���{ऌ�6�!�$���68b���Y���;F��5�!�č�k"��o�	�bö�+9k!��	���P3���K��X3��BB!�D�!v�y�e��Y�tۄ.Ɵ�!򄎓OT���ی;� ����x��In2�"<E�d+[7#�j���ҵD�|h�Vc�y�bЏP%�	pS)�lD���� �Ԙ'E����՞DISj�1mdF"�׳=���=��'���a�l%}�YJ�!ú!�"L�	�'Z�eY*�0h|8if\92���dV���I'�p�B*�o4����Ԗ&���U�d
2�`ǥ�+]u��Bbo��A@�
Ox�`!LS�$���B��$����t�'W\|��y�㏃m�A�WoSo�.$��j޴�!𤛼J�f����W��h�>�a{b���6V�`���K�S	h��m��
�!�dԣP6�p�8K�reS�(�E��O?A�d��`N�2���1-��*��f�<���6"_\m�"BD�Y������b~re��0>��.ެ&��'���g|�� #��Z�<	���Y�(M�A���}IഇEY�<yUo�%c���늉bPȕ.UX��p�e�$�I�W埠D�
�#E�<'C��$[�H	l���ݑ�*�U����BM'�S��6OL9���.)�0�hg�0_���`"O�lʐ�ʝ@���A33�b�$ɍf�'�&�	�U�'9P������\s*Ys�ܬ��D'�S�2�<���ĚO�������S���䓺K�M�,ONO�gy"�ũo�~T≍�R'<i���Ê�HOT➘��E+?�PF�r�H=X��W> 5�9q� d�'4a{)�9Kl�R���D�*H�q,I*�M;ߴ��O�'���1Iخ���&�*+?l�j�.����	(��$0�P�r�/6o)f��-�!�����Y�'��,:�/ވ�4m1��#.��B��$Z��0|�!��ӀD��-F1:L�AՀ�A?�J̦Gy�&�	F}0�  ���`Ǫ�X�����7�OF?�yJ?Q����g���Ѹi�څ�S U:��Y��Mh����}B�'�D}A�g��-���2��i� xX.O��h�&lx��ԖxB�O�t��㟼 H!�Z8,>�����#%~,��׋-�x2�Z�0�P��oɌR0ݑ�@#��	+��@}���eS��?!�Z��'%2L�g~�U'Cvm��+�
".�J�����<���W&��'��\�I���e�]�f�a�^�Ze&�D�E%�9�'�ؖ��'��'�dRg��J���3&����� +��_}�:*��]Rp%ޟ3���`u�� ^>��BO��`����e��z��k6cW�`Ұ�=���'
d4)U��6'�&&�͒@� ��RTy[��cA�8a�OX pi%�7%�"ꧠ�� �a�$xHX��* �=v��"O�4k�C�m�F�H�j]��@ 
��.(���t�N��5��
G��6q&V�CEbEo�$��e(�Y��+���ۧ]�a}"`ͶK��M#̃4{@!�� �Ix����׽'dQ��U t���4g�,K�t�c2a6O�R��S���ʡ,�=9P�BG鉺X�B�
'���L�p����&n��UhT+t\��[%C���Tls�G�8�5��%\?�xb,ƢjCrA ceX`��9ppH�9J�`$�Fd�5Z��Q&�^�B�Ӕ��!oIb]#[���,e�
ղav�-	׋�;ZP� "O
��#��!|&�#�^6U�d�%�;�X�C�4��Y+�'Z���Z�#z(�s�J_5��I�%{�ϐ��2I����W�d��Ҏn�<�k]�8��(��	Jݚ����6��+��Q���`�.,�����?�p<!S�ޔ8r��g�H7�
��f�'�r<��&�/}4���o��|$¥ꆐIlɳ��I��0c��r��Ă�Ew-�=��-�@ �E�M� Z����)I��Ò턠]���j%X�x��|�p��?(�R �%LM.!X��y7�V ��a�¤(�@h&
$�y⪝�E��$��$��������t��:KB]8���[HA���O��8�ӄ�"��ӼӃ ٬�JmX�(�)u�n�ȅ�QB��#�,I�����xjtť y0�S%�W��Й ���E�^@2�Ǔ<Ww~��Qˁ��O���-����B��;\��y'��0�8ɣ�I� |8EC�eV�s����LN�+dPe0��4Yl�C[ &���Jk�`�p"/ӞS5�Q(2����	�N~�P�,O<d"AJ޺d��t�%G�70����&��c��K^s�xÊ܀x�4tq*^:d��O���`��
QB�QS$(Z;����)F(o�	��ڴF����ד1��0Te�5Y����W�X�!x±�0CލBV�7��<���'�l�����X���k�,N9�J\�1�F-B�x�ѓ��)#��@yu��,H0DB䉮ޢy��JA[�Р�g㎑Zu�6��4M>R9�Q�[5�b�Q�+�[#�m�������%>��<CÖٸpEa~��BU4�����V�����Y��sNC�����}��U�S�,��n��A������;i�H9�1<∜�{���!T��#բY�x�(�$['��O�J��S+�E���3RE�]B*� U��p��E]ޒ���2K�^d�`�	B�Dԁ%��Xf)��I!�,%�1lx6�R	i�7M]�~2�e�(��f��#�"We7|P@���l�⑎�0]Ez!���S"?^���QYJ�B�ɷ[�f�#�_Iv\�kjX�ؚ|�e�֋6��=�$�U�G���j��	6X�j�3��&�y]w���R�-i��#V̉)f�r��3�Ѱ�4񙆯2�O�m�#-%xĂ%A�*�qo���A�^0KT�@R"!�F�3�fL	�5�4��
%$5:"��qm�ԡ��$Ex?*H� '�#��A��e�ay���%@r1x��!	��C���rI[�1#�l
��Π�T6��.hI�"F���=�G�@+(C�A�B�V�nǤ�h��D~R�J�՜Q�ш�:�&Pe�ȺhT�b?��m��(��`���۳M����=�O�Ԕ'�|�!��G�x�f��Ϋ����)�� =p��+�q��a��2�$�Hc@G��	#?Q�JO���i���D	^4��b̓_6�$�l��`�Z0�ɊT{����ЊA�R��U�f�X�Q.�MCa�C"mUؑ��O��dC�yX�1wCLk>呲Bܡq�'��h�S�E�@�hlZxo��&?YH��џ2���np�eI��I?:85
6�'!���Y�z�Z�@��SO�8;��l�e�W-��P0�Q�6r�'�&H0�w�0h���R��!�X
y�����'.2�)Ip�ц��<�9�䟡t���ꔠ��m����ßb'/*L��?�ɨX�&,��	=(]&��F�}5h���yZ�p�g��7�h���Kt$�b���sn��A��A:
g����'NX�(ǖxr�I�kS@��m�v/�`"nT���OZ`��ݫ-�����(��e���%�c��
4H<`�Q��j���Ii���	�bK���*���$V0=�����t,�,lZ�_�l���C�D��\�|�Īg~Ƙ�l��̃�ߤx�v�k�M���xro[�_��1���C�Q�)��s'4%ʵ(�x[�9! �v��4'b�'��	����Mw	�~Y���Y+'��4�M�H�<4K��� 2�!"2�߶ ��	$�#?
����ޣWP40Z�I�zۆ �M[K)�d�<R@�l.��U���1rM����.��H�����`&6���R/�>RO4��s���k�Դ2"L41�x��5oZ?��fgݸ�Y��%}Zw��j�ڧƑ�%�vh��n	�ly�p�'�tʓ��D��i0fAc�.�";�9�����@��'t�1#�2"���O"yɇ�KqF �D쑭}��$b��'y�I�G��	~�'w�.Y�'�q�����]�t���*Fg�(���*w͟�K�A@�r���#��A�b@��Zg��X!�'�o�i?A��'������0#�J��(�ǺK�OC��[���_B��G0�<���0қ�;O� b$����$P��q��BŢY����#)�ybO�))^<��랯;�`�OVq�������oa��Z�A@	[2~�[Q���'�q�l0E��f�>���D�2?�QV�O�4[�'%����gȲ��Ϙ'\������D�f�s�mJ^/2�
�'_~��	��9�D���H��Md��*�'_
�s�'?�4��B�uS8h1��$;<�,�1�������v۪,UZ N���yr-�{���!�`��{.Z)���~����c��|��
������*Ȁ,�'�٩R�~]�!"O�=!K�_J>T����;Kz���x�V��>q����'�l	�0�Y�S�j�kr��u���;�Ԩ��A(#�e�Ta��&Þ�X�B ,H�r�~�(��	�l�21�D��$A@�)Ge5:G|���'R�x �$�<᤟HiX�$�n�������k�0t�b"O؉bK��c�Y��IZ�_m6E�ӎ�8!�`<���Y�N��1��FĦ�G��3��M+�@G����C��P���l���Ʌ�x��bT�W�� �	O��6��_���`��Z?����VfҴ�I���)p���dcQ��C&��d	ڤ�	-�����gkx7)C�a����ƴs�����3N_�|;:OnH3w�'� �'ߓ5&�aC��F�^]�=�1�v��Ta��<���!Qܟ�re5��["DP�6��u���n�Hh�C"Oj$ӣ�-�	�NXa�[j�Oj�D�!v����Mۉ�	��i��|�I�>�<��(8&!�$�%�9)���z|B�`u�� ��+S?��1�U����?c��!�
؝�޴C0d�A��z�d1D��)�$�
�Lm��˭J��q�qB,���-J����Ӣmft�1AN�=*:�1�c��vR�2���mg̲1�ұ\P]8`[�;��,��'���"�OnL�#�îl�$�"M�Xm��ú�>3:�?��'�`�q}d�t\�� Qd�M�r��4�7�0=!"�"�	�-d��g��a�!�Uo\9O5O��	��?!���W=B��99�'��~�1؆(�:�ў�Gy򣮟��P�H�6=A�j�?&��$ ��^��?��OV�S�g≯]��� 3��'W$V���=M֘b��Er�'��H����	#/V�
C�G�[���MN��' x�b"K�&}�Ui�)O,پ�s��>��*��l���M{����8�WB�MSc87�|[q�'����$�-Q�@��-[9�,�7bހP���F��������2m9�i��)�*9"0���!m�PR��a��㘯K4P�EŢaH���Ab/�M�e9O�O�g�;��h㇀p�^8��bP�3���6
��d�� �BZ(:�r0��A?T�Y�I,?)6�'�2���b�g�RTo%]
�  J���N>	�{�^>�#S�/]e��@48 ��!&�O<�ɓOJ��6�S�N�䕂�C!oenB�ɛ^�`��ű����� �p� B�	�Ts���H� z�j�p��LB��8XF�c�NǞytsӈˊI�*B�ɍD�򙂴��
o,�E;�@ܙq��B��'L��PJ��g��AS��	��C䉨{7�-���S0@Uk!M�'-6�B䉫p�΁�4�\�H=c6�F-6��B��y���j��6;,ڐ�D�sfB�I3FJ��C�c�Eo�\��^�_�B䉪s��A�B�{���#F���.{��?Q�+�'7�j�t��{�:5� l�FH��ȓX��Ƀ%!�w(� ruBΪo����'�R�	��>16/6ڧ%�ޡ�bɝ?2���קN�8��ȓ]�v���D�w������_�4 �'!h!�����4NT�r��M/Y� lQ�E�XC���D˺7)��2DF�'�H�0��$�ȑ��Bǣ	�LKǩDHH<Qփ��t�X��l�hcX�{���^�<��m���+��� �vn�C�<1��û ��S��(`U�d
��y�<� �J"h@02�J�q�jȡe����5"OD ��I8\v��aoV�c��W"On��4�ܮ$��5)����[|���"O&D�fԖ3dPW ��fl�$�"O�UZt;q�.�3W�]N�"g"O���5i��h�,�A�@�>_��X"O���~��ؑ ���54Af"Ot���b�s�hy��I�>T9�"O�l	aȗ!QX�H��w����'"Ob�R���2B��Hӧ
�q����P"O�9Ze���X�vS�I��'"O��aVa]�I��ܩ`�ʯx�9sP"OԸ�֋=o����ԗG2D�"O:���d��N�&����$S�X)�"O8�5J8N� [�J_�.�4z3"O Kd�_FE6�A	����t��"O�q 	�&{A(�iվZ{�(�"O����m�"���b4HC�[X��g"O�uzSd٨.�~ڶ��P�FH��"O6 �&��#���$��\NDpQ"O�HzBO;hO|����6X�H�v"O.�����e,�$C�I�6l�~��r"O!��� �J)(H�;S�B�g"O6U�s	�Z٤�A�M�b�J}Y�"O� �@9ZﰽR�gR1Z� 5"O<�i�.�k>zY�G�u��aX4"O~h� 'ߧWz��ֆ�N���"Ol�������Lq��tj�$ٗ"O�I�� QN��x����0X�+�"O�,Y3eJ��PH2 W Kf%(t"O<\YRf�	8,�Y��މ]��)�"O��sŊ�v��ep�n��A�໠"O<�q` ��h	bB�,�"�%"O
��Bl�* ����&�#,�:�C�"O��� �/�聥��6W@�[C"O�w�1M�q������"Oh�	W Pd�q����lQp�"O<%q6�͕~q����LyP�"O|�r*��x�~����98�\(�"O��#�A�@�ʱB�mÄbxh�[`"OZ�KD�
L��ʕ��tSz�A2"O�HY�l[LTx��5�D�E��i�"O�����?��t`u��	\�8Ȓ"ObY󀡁�]d�q�ȕ�YE�9�s"O���Gk�2.ƖD hN,
Q����"O�g@Q{fys�	�o&jŃV"O2m�J�.7|>5#$	C/.D%hq"O�\3C�1j�2k�	�
Z�%"O�EC�"d:�H&G�R<�M�2"O��1�ӣl���4��� ��"O�xa�$J; ~V���G�$��"O��PkĆ���&�,3�JjB"O0�Q!�:{�`����Şa��Tۗ"O� ��D�|�&�r��>X�� xQ"O وE�J:z\m��,1 �X�"OZ��So�%��*��ͧ,3v�"O&񛵫��]dB1��&�e�� "Oz�)��[�q�UHSě,�:0v"Opt�d�!8��з惴7r,SR"O蝨5F�&dz�O,GL��p"Od�����v�d1�'�5(#$E �"OZ-���`�hPv@U�}�.|@��B�<	F̀6`;���! N?������}�<YWJL�>|t�i���2y��c���B�<� �	 KCh�$X1BA�h�X��S"O�Ȑ�����+��B�7�X����	���B��'�P�0��ALp�90�ZM��Ch=�d)�^��T�_%�d����N�X��@AEO4�S�O��Y[��0-	��S��2:�,A�"O>�3�ڃ3.�0qЁ�n�|Y�W��a�EI;`lsp��b8��H`��/'�����/�,y|�ᰍ �O��B!��X�;�b��zd�F2P>yc5 û0)�Cቺ���`�ݾH�Fik��[�Ɇ#=Yf��KWP4�u��ǸO_� c���D��@e�dY��'?�qz4�3z		�u�ޡ�n!��'EĤ�W���Y��֧���eV�T��e��,c�zx:�Y=�y�i�5]ڈ(�d�;j	Ԥ��G9�y��ȣMa��V�L�n{n���ɂC�Z�j�14#���1�ܸvb��Ğ�B�ҽ�#@#U�V��5K�J	R�Cw� π�ɀ�E��Px'��}bU�u��@�
��OT5���O?E��8��K
���O�~Ȣ�T:��� Jh���'�P5��R8�� ��HN9��ꕯ�"z�2e��.Α~���S��y�#��PVH�7�ˠE����A.��y��GL��8��K_�:���#	��y"KL2~��u��L :��y)^�;���X��>��3�Q��0>��	ܝ4�<єo�Z�ș�� �=���Њ��Y�����{�
J,GF��"f��~�O?�`����Cp~5JA/ tґˋ�κppt�0��V���?y���:$xܔuiI1{� ᔥMU���k�G���Ӗ�(��pM�ݒ��K$���&k��	�䙬[��P20 !}���'�r�zV��#F��e�w�E!�h� mǩd�$%RT˞'|X��I0S⢕)R_�+t �8���2;��
�T�#�G�y2o)p��mZ�(p�x"�C71�.�@�v�zsÕ�V�j���2��C�I'Y:���+��v���Ǌ�1,��7�'u�rp����0�VRF���H�\J'�7�s��sr���* 89�⍘p�,�0�=D���ԥKQ��ʵ��'e0ܫ��߯@Tm��Eʮ]^�(Qr&C=hx��sQ���W�OWj�P�m� RU�XӴ$�>Z��e��I�"�x��6�R�-F�2�j�K���p�
�)�@�3)ĮP�~-���ȟͤ��
� ӕ� e2xɢ�RnلPFy���$0��N d6t��SkӐpR � 0Y:TH@�C�}6(�V�R�W#���?�TБ��[� �!Qv��&����<��uXϑ�e%�!0�<�Zȹ��;���Y�C�ܻ �TP��Cܐ-�D��$"Ov@��ܢ^��$$,��0�F�G?��1��P�MN�l��(I�j��).b��b����J�)�47ᑔ'7
�yB*�|8��4戫M��XPI�6	$�4i���"��#�ʛ6�d]<Ka��^ �{"�ӛ3����&+'�d4��Ϡ�(O��EF0����i���}ђ-E�F(M.H1!��+�*`��*R�0M
��ǻ53�y��"P� C *M>���*���Mc�ěO#|�P�eӻlR�põI�ax��@�œ:nV�t�'J���w���Թ���ڼ����+O.�C�j���=Q2
 � h��"�%�I r�WY�	�9F �p$��3K�?%{eI6D��
�`#3B����+D��b�V�q���B�dѸ��)@d��O2$��a�e�g��O*Zq�thL�`p5x0���*�C�	
Tw���^.o���;� gV�yǋ94�����'��Y����)ؓ�֕U�Z��k8��3@�/(��˓7��Ѐc��Ԅ�&�x�ن�,(6%JTEM�v� M!�F3�T=&��2��-j�R��'�����Z`ܧ(P��	}�@��������������K�9M�n��K�
b����p/M,�M3�I�rip!lR���O^�)L�:���A? ��b�J�o�֭�ē��0�%���oJ���P�]�<���Ү��_�V�І�J�'Ѝ�3,ߑ*�Ȣ?�p��01z�9q$��/�y+%�Lrx�<adO
-�}o��f��J�[�.�vP)4H�_8$���_6g��-ʢ�'�v�#7�ے�x�ㄳe3l �y���d1h$�ɻp��� 
U9�O�.�w!΋��Q�QQ��L�'m:�FT.�0yG�H� ��Ov5�p�n2�PbH�"}����2Ku��@��x����WlZy�<q�ɂ��QDiS�I��S�'�/��I&<�4AgD����g�S�? �����J�)e��B��JU��u���'�pe�!�
}� 53����r�X��rbU�B?������s���	�IV���!#�P62�l
֍:�N���h%�Q������,�dT�l=L �5er�	S"O�X�p �>i���B�FW�tl��#�W��맪I�_ֵ%��|Z���T��`�H�����ƥM�<4��
+�ܸ�+1�f ����C̓�b���:Or�9���X���f�?QP���"OJԛ�"� N�� #�
K!}ĸ 7"O���%_����V)��8n4ܚ���-/�v%8����]/P!S��
8�轑�F-<!�D���`�K�vqn1I1D��.7�$�*]x��S�)��ӡt���p	�s�.�R��%2odC���dJq��%l��h	jG|UF�K���b�T �����ޣ��2!��$�NDJ��� Y�a~�� -V�
����eQ2mؐ��54��� Ɇ�{�6y�*��JU���b��׀X�O� G|r�йE��M�`�lܧT��t��z��(I�Rj�D݆�$m����+�+6�D�0U���V)�;�̑S�U�P�Jӧ����x����{b�h�`"T"O�9�D�Y2* �THq�L!(�H�`���`��E�D\�����'� h׍�T̊-J�ʆ)/h&�	�5¤�� ں%�
Ԡw�T��&
�)v���CRbO^��D�� FxQ@ʶsbt�dA5Bm�̃@� �l&\�f���x׶�P�^.���b�ڻ)�!�$��jD�i6�$z_���5h���γ�*���-��ӠA%��bQ/�<�z<Y�'��Eh�B�I 
h9$"��p= l�"˙5a�6Ox�����<9#���,�R	jӪ�;�$���CK�<���2D:����6`�L�J�B}�<i�eq��*�g��Cʹ�
&��!򄚄*,R�A��O�g�|�@T׵J�!�D�!j�*��Ŗ!K-8�&�l�!�ȷQ�	�'$�>K1�+f�_2!��6�Ph�Ʌ�,u���S6R�!�[~��5�U��BU0B�(�!��	Jx$r����k��5#�@�1!���U� ��B�è9�m7O,L�!�$R�er^,����6=�B(�4���|m!��D&
@f���Eڬ	k�\�$��7m!�d\�&�v�yV/C�/fV8��>ZM!�Aj*��1PÜ�SP�l�I6�!���3A���#ɕ9�n1C�&�6�!�d�d6�ؔ�V"u�򝁔.�=�!򄌩A�������\�SJW#�!�$O�C�Ft 1MO����']9�!�x0J@	,���b��}�!�f��3��s�L	�VB��Q�!򤚔V��x���'a�lт��+�!�DK��.Ku��7,��IJR�5�!�D�o+����<9�
���̓z!��߶Ro�2�ŀ�vÞ��
��d�!��� ����7�bU٣���!򄖔g,dp��U�@0� '��[l!�d@1>��y�Ä:BY�P�#ϦfH!�̒w��5"����:4Jxؔ�ҔV#!�4e�z�	U����t��B\�!�E���+�88�ԣk�O�!�<8 N5(�(�l��`
v�!����E��+�!����*Ĳ0�!��T@��]Ej��zL�$�D.�|�!�<4���і;7|T3$��^�!�D�8}:���E˖-8��!P	e!���1(���b�m
�)�d�k�E	�Ik!�� ��C0�!n��2��TغỀ"O�{#c�d��5�Β�"O�9��l\6��8!�ԙ_�0�P "O"�HF@&&o���b�e��xҦ"O��q�Ӥ	Y,i�Pc����E"O�U�:p�!W�%
'�4h}!�ɖ.φ��k�1FsAJ�/V!�����,�Q*֚uƬ�V�4G_!�Đ�{І�#+��WТ,��*V!��y��eQ�6`$	Z�
Z�%V!��ϧy��Q[�G�T9�5�E���=/!���9^�E�'B��(�*��`�!�dJ+e���P"�N�l7p�"*@�.�!�d>Ud����z)�@W T�!�ۅZ�8���fٲ%��酯�7S�!�JVyZ�"Q�W�2Dq��^�G�!��A�&��	�=�b-��,��b!��[
B���*1芻V�z우�ψ6e!��� AM`��u�:b� ��C��!�DM�Sd6����*MD��TAЛy�!�D،Y,3���h.�[3C�-�����>a`��˾l�Ԍ/�>�Ѩ-��(1��?�l�@P\}�o	a�B��w�ǀZ��Oq�����UQ���5�հk9 y�W��z�'�W¬�H<��M#�O��0tL��n�p��,T"l���'�°0�Ȇ��M��'~a�TK��[T
�r�ѶP�2���j�4�&�U���1���?A+��<�'�$��';�ݘ�
��%�X�'>^�X�!�I���u��Y���K���i�R��~�$�ÈKW,x�V��fh��@�7MC8��d�<���I�a�t����j0�/Τ�1d���$�'C�<����7;F��N|nZ�I� ��D�I��[T�D�Vu2�rN>LRgO�"& ����OR���MFh,0�dX�$.a(��,��`�q���sK��秨�XPrQJ�nb���,�4IT�E(��E���T�F ֩��$%�Ӥ*� ��_Jbs̖&{��!�A��_�HP�ѡ6�nm��5���DE�Sr��'��90̥B�Ҝh�"	�iH<"����?!�
�	f.�d��6O�?�+��Y�s���6	æ;K�l���O�12Gʝ�o�2h&��~��J����#�K��p�8x'����`�q�[�������E�4\?-�$Cea��3h��29R�j��I36d�'�����ѪV�a���\$d�A�	��)i�N^�i:�IOqB�0l	v�PI�'G�Q>QB1����专���L�T�5��O�I!�;�
ô5Y"آ�"M�~ɦ`@d�R��Gc�:�Ɯ�LJ�DG,��� ���<�� ޠ`����Vg^4 ����}�	(٪~kb!x.O?���A">%�i�# L��0���uw*�4��^��<
Є����C�Oq��&A\�f�l0��� :���R'X�i�1`�'ҵP���J>Y��/�*�:	*��ձtF*H���%?���	9\���;Ba��iUO�OLm�Q�h��s�Ù�(��YЄq��0�� �p/t<�D Ř>
�?i�R(T�H�����F�=�P"�)��M#��=8�� �ǒ���S�����+]�T�V������ ڈC��-��,���ƺ}wD@���h��B䉨s�=����tM��$-��$�DC�{�L���Q� ��cO>$h,C� L	��'´K >��&,�"�>C�I�~��$Q��D�m`�h�Jb�C��$z������F h"��K��ƙd�C��9O8�N�^�ք@N@X�C�ɩ;k�p�"E*ؘTD��5��C�I�@�6�pg(Oz�h�H��bĨC�I1S�j�#Uj�~�^أE�܇gw�B䉃A,QH�DǪ4�,|+�W�=��B�	:rT����l��-Ӹ<Z�mR l��d��Ta2�3㎣v=����	+_�!�d�vbT�c�a�!T9�Y!FȖ�YW!�d(j�A�N?#���1�Ȍyo!�Һ7�YƯ!�V9`o� Jx!�$�$�^���Hdvl1���ۘY!�d
��ҘkG�,nq\hb��ʀ�!�� ��蕁W�JL�\jW�:��A2�"Ot����ܸA���15�;bJ�uC`"O>�"�M	�($�qġM=9a�"O���R8'8�tK��[����B�"O2���D\���<P���*:��x��"ONXJ@�F?Z���"f�Ө0�1"O�QWn��C`�vg�$���"O��Q��+:�}��?���"Orr���$T"�RRN�(h6�r2"O�< �+16أ��7����"OP�s��mH1BW̍犙�gIV�<I� F;J�B����"`�<�3�UR�<a�+�#2BQ���
?4U"�h�<�N��tX ���`�P+Vh�<Y�]�1�f� ���(j&Ud`}�<Y�h�
*�����P�l�P�[w�<��ƕZ�eA��I?t������s�<���8-o������;v�ڝ���q�<i2	�0Zp�Ƙ�r2E2��C�<�%��8	��x�E�u%�6[}�<�āY��9��Oi
� v�~�<��˙"M ��F*X�z% VJv�<�vϵe4�Y�$i�='J `p�l�<	�D�4���\�}����F�e�<���0{�:�p�-?�v����c�<IC/1�^d��`�^�؋�g�V�<���_]EBP��(����Qx�.�P�<����!KH���h�NػEv�<�P
�&t`��8TJ��/l��;u�o�<9f��0g��@r�q��K�hRk�<�󠂡*T�qqa)�o��PP��Q�<����H��$�?;p	�G
�h�<�%�_�b �Noer�;Á�e�<�PCE�.8�T97F�;���j�I�<yg�6�d*"M�����fVF�<�T&�t���JFU�N�Y*4��A�<qF�÷F����/�'w��9���<	 b�1r��3D�q2��}�<���W�֭�mG�,m ��y�<ia�[������t
���D�Lx�<�F ��hk4M =��sԂ\p�<��b��S,�t�7�"<x��KbK�W�<��K� �Ɖ���F4 ���� m�<q0��.(�h"��_�1�2I�wJh�<1�����.=�uA׀
����^|�<Atm��J���3I٢J�X		$�VT�<)@
+p�8����`0����C�N�<tJM�8����L[�4@�G�<i hm��]h ��=<#��;R"�A�<�p,MM�Z,��A��Xډ�
�@�<y�H=4tU#s�T7s^YӶ��E�<��Mա9��
�0t,�eQ � @�<Y��T9|�p����ܕj}����FU�<�^�����\ R�8�'�A[����Y�ʉ��G���@�͜>LD��+���]�$ٮ��f�B8F���T^�!�2`�]�(ĳR,\�*T>�ȓ ܸ`���N�����KG15>h��wf��D�1W��q矬\1��)�x�r�eҞ �[6�*��ȓ-�pl;���,N9�=�%%��R�a�ȓ`���@��|¨��Se�_(x��N4�-�э؛���"�� E�B�ɭcIA�#��2I6���Ua�)��B�)� (y�጑�$;E;�N��L�*V"OH]sOA �Q`-�,֎u�7"O|)m����58�����h�"O���C
"�>
�#E�`�T"OP�q$n�+��,8��v��	b�"O��zC�!w�Pa�7A��q� �V"O0���dR��je�S:) X�T"Otm��ʟ*,�CS��=L�N4�"O0(S5�ۡ$i�ܚ�ǝBl���"O���	��؜@r����)h�"O���A��&4�0  F����a��"O�}�bC�� C6��<6<(x3`"OT[ꉋ-34�8�#C(�2"O��0 D�N�
Q3�T�M-(��"O���`ǻU:��hWᕌ�B��q"O�����_�yK��+U`��thc""OD���^�<�JO�c8���"OLJ�A�4^��D�2� �>ԅ��"O(�Jp�T�b��Ul�>��p"Od=�奝�Cjv�(ӋE9>!����"O0d�V9���Ž0��h"O&�eA��96�(g�"G���"O�-ӆ�K"�,z�lхE���"OF$�Gq�1�bU0�~a( "O�D�c�^�s~pH���ț?,Z��4"Oʠ�'������!�=��*"O��ag�_"y/Ƒa��2}j�"O.m�t�R��d������Pb���"O11�)ѭ�����uU�ՠ "O�Q�Z'_yDK*X�T82�2"O|P��ߡ,���bi��6�r�"O2��ba� `8H��!&Q:XN� ""ONe�7oDC�h܊�E 5"E2�"O�<R�	�@�(�$�'%��Y�"O��� H�#G�X��%��|J��`"O�!#B叇������g�~���"Oځ��FThi���ĭ��	.����"Ot�a�͜�%眖.8����B^>�y��Nn�	�IG�7�ʴb���yr	�`-��#���5ŰıE���y�#F>~�bp�'d�#en���'��y�,��q� wϮ[��U�V���yϧ &�����V�QDP��A���y"/�nC�H8͕�U�8Ӏh�"�yb��Y��H2d�L/h����Y��y�HQ׸�c4	HF��DX��>�y��V+0`����Ʊ�vŠ#h��y�,�49� Dd ���Ks,���y2!ܞ=��]��&I�}Q������y2�  4���#��;q�nY�
�y2ƈU�|�0�j�2i#E���y��K��;�L�N;\�̕�yB��8>�����R�s��9�ӡA3�y �&��mR�@�q8���Ց�y"�5�N�@��P�p(�T��y���'i����Cj�e������y®��.6�0�t��^+����?�yrG@�N|Ik��F:�M'�J(�yr��NBB��w.�P��Mr���0�y�B�� 5��a��E��L���L�y���(q�|�:�FJ�D����&��y�GO��p��ʡ=˘u�Lɭ�y�kT#[&e;dD�7�h�qc+��y�(�R�v|!�DU�*�~eb���y
� �� ��3k�)A�>�M�d"OTy�w��n)�5�&"յA���Д"O�p��	VSД�T�[�hG���s"O^ȂB�A�s�\�gȕ'w/�a��"O^0C�)�_wDl(���;5>��Q"O䌓��H������i�9�"O�T�s"L�nwtx�bć��晨�"Of,�$��ps�8��I^�m���ip"OF�a'E�"R�i�͟
LFt�c"OT`bG��UP��;�F���\1R"O|��a
�?P�]h$�K����u"O$	A$�S��,Z��@��$;e"O\\p0E̶!ujq�R�[�T�"�"O~�ʥ)�rE���딶 �,�H"O�2�n�/����G	���i�"Op��ȗ18� Sq͖�G'z�x�*O<�*�5-=�4&iF�����'v���Y4*� !�`
J�V��'�Zt9T��P�l0��C14u4!��'����� X�b�Z(`�.`U���'n���?1+�a�쉉D���'��Ԡҭ'7
��5��16޲X�
�'0>�n(%2*jU�ֿ]�*��	�'��r#�x�0Q��MW �|��	�'
�͛7��y��`����Z����'$�u�!c�
�TIg$�~< ��'l��`��o��бj�<Ɣ�'H�v'ȧP^����nH��
pB�'�TlccmѴj���z�i���y�
�'��]����<N��1!������R
�'rܨ�2�6f������;����	�'�F}�Cƴ>�T0��Ć����'��%�S��x�7J�8p� �{�'X�B&a�w��$�7��5���b�'�t�b���-M��#F���
%y��'�2�H#�\��0�+f�C�����'�>�QWpf���VA�0�
�'Q�Xh!lӲ'0�q�v%.D��
�'�K[%/�(&�tf�)q.�N�<6��s��+��;V�Դ9�)VU�<���ӎ_N���fK2NcldA��HF�<��ȋ�,2-xbձ^<��p
I�<q��˧�0�r�bSF����5��A�<1��
8�p����Y��Ԩ���c�<�"'�)&�.P3v�O}>0;uEi�<��g�'	&�� �뗩?t � &i�<Y7�ˑK9l�P�+�(DW��B�E9T��F"="Е.�������0D����D�%X�<&��Z��1D�h�r���&K���L�.�00n	����Opã��@t�?�U Ѕ.��d��D��,8X�E	жq�V�C�<��и��[�k�.���Pwϊ-Z!�#�m}"Ê&Iv�I�1$���$���c��9�Jq �_�% �m")O�J��'כƞ~���l��禁)�]08�� �G�(���S��54��4h�-\�yI�f�
(��-������y2j]�x�D61��O+����<A�#�f�X��5O�$�K��2a�$e�� ��'�JL �����y��'1d�0A��5�a�N�&:a�	����>l��H!H7�O8�"���X_n�
��ݻk&d]BO8L���3 Tmreb�>��?����צuZǫ	�s�uu���n&R%��V��?yкi��]�D�ID��?�1��ԌW�`��V�˰2(DY��J!}��I��'�H�a�	�$4�n�C˝C�ԉ�J� ��+^�M+O��X�JIF���>��J�r�� p�)%Ӟ�9̎S?1���+�Hϓ�?qe��!M��Be��+/��s�����E	",�P�'/���&Ǒ+oY�ID��	q�T4���X�R5�����J)7NQ�E��u�����3}z��'(�6M�O��=� �Enńk���B�Y�20�A�O|��<�+O�>��ĊH�d(�`9b�0W ����<��J��u�2O �롿i�|micH����F�������]��?ё�i�yQ�b��[���ӷ@#6u�'� A{BV�l��x�%�?D�$�X�,�Ob��e�J�T�h�xF=O���^�
1[J�|hW��<�dHa�eP9W"SaD�>9��+��1f���6�C�(�ԍ�4`��#$�p�Ǧ��9��ЛS�)���O�����	|�O��F٫ I�!#kۏ=Q��O�D��p���'�,�͊32,�e�Cڔ����o��K����MH>��N5!�e�*^�j�@��	mD��ϓ��ݏ\�-*0�%��<n���h���#*�0�E'j�|��բ ���	ɟp:�)
�`<�y��0�����q���( PU!�&�4c�ʩ����q�R$ђ_f��K嫘c��>�>O�3�Oԭ�4E��L/u���hM5�M���k!0 ����?���Iɟto�� ��@!G�ΜZ�h����L�&�N)(���s���+u�TC�,��g��(1��C�S�<���ǟh5�6�|B��4���HyB�2��R�K��YD�Z��eWv��m�7G��O�Y�v�W�-X��O��Kp�\�g����s� �2���Ӊ%��Ұ�͟��ȇ�47�D CB�l�D��D�լZ}9�ŗ�P�X��ʙy�S��;O�Ҧ�i�R�pW%N	�<�:��/\T�
�/�O�%� ��ߟ�%���OTVh���4l����RBl!
ϓ#��O�T�)��� ������PnB���*+hd�$;��{�"���x}2�ۘ+ d  �=^���2|@ii�e��Od\a��@̴QB�� D��>�t��]A�6W�������u��'E�ɔ*&�Ar��1���k7�F���E�P�Y�am���	�:��]2����OI�	SCß���%���|�L����!: ����P�!��5��DN?/x��q%�,3>���4i+(�J%�C��y�'�d�@���?�a�i�2��q�E�[��J�$�&8�q�O��D3�)�R}2eY�Z�����gIC��Y#�
��>}���'TUhDZ�V*�x�-��O��xa��0U)���.Oʬp��հ�~b���/M����5TA��Ͳ@�<�Z.��R��4��"dFпez���S�do �� ��҅�P�A���S��>t	 ��䴓&nB
j5J��m��!��ny�i9�5�gj�w�j���Nݕ�p��'�ؚ��?��i8��3� 体��^�X��D�0�A2E�{y��'��)�?�ՂܐP������C�m�}[&k�Y���l�I7
�����O
xoZ��p<43@U��Ͳ�L]�C\�x.�O��'��]q@a���O���4�
�pA�E���=[Dm�@Ǹ�gg�P��3l��}`w��&�p<!��'�T��
 6r��}Z&hZ�05��3R���R�
4�S�u�N}'>�=���	���f�^�Ilv��g�7:N�6�O8�#'��O���~�'�"�im�XB�gFD<�֠��Jٻ�{�',D�K�2��R&��0����v�������MsN>���-Oh�:��{�M
F�R�Ix�Y���(E��	���9��!�u�L��y��'��;d���%�E5&*8� ☗JL�1cL�,�p>�� �2�,> 5xB��2z��� ��Ӕ0B��_V��j�jƓ&]�#>��Qئ��aƞ0��i��f�As֠��ȏ�?���i1RX���IZ��?���Οf]�M��쁻?Ǟ�T���$G}�#��E�z��0b��y(y�QH�#I~�'6F��1�' �@!� `�U��O}�N�A'�!Ã�q����G��~�G6�d}۟'���='1�a��o$v���O��5��j��Vȭ(�Gݨb�"m�����l�XP�S*"�F�2-E�N���2b�v��ªŢt�v�$
5;&���o�O���`���\�F`Q�Y01�ĵ�cCT{�:u��Ɵ|'��G��č�\Cn��eٹҘ���a��������ZXH��4���F�Ng�l� �-p ! љ|2�iI���4�3?���4 "  ��|Jd�Z����5��O�d�^���h�Iy�I!������ c� ӆ�]Y�%!�
�	��F� �O��u��5��HвY�"8R����Z!�9�����M�;R�p� @�?�'���wk�՛@ ��Z,}�ⵆȓ���J�j�0E�a��MV�0�(}�ȓL������D�QO��[e�6�(��ȓ@NT�6��:P2�O�%H���S�? \��� E~����$pV�l��"O6�����	6�칹W��+Bl��V"O����n?(��YTD��_@�4Q�"O�5�я���E��"ߩ�pЉ"OF���+9�\Q#^2C&� +"O�q�S��S�Ҡq��=(���"O:ܠg'�:@)\�`%\:1[VQ�"O�  "�- !� �@�����&"O�zG\-*O:�j� �u�JI�"O� �P-�+�0E;�Γ{ն8�"OD�P6�M��I$i�1�'"O��0���
����mW*lHIP�"O��Bug_�}9�s��)njRld"O����A)$��xaN�zm���"O��Aa��!L'�2�N=kXi!�"O��ذ/�3j��)�X�1a���C"O�Sul�J09v��$i�i�"O�e2���*^ S� �
?���G"O�i#� Ί8��'���<�D|��"O H��]�U����n����"OR���:f��\z̌|���0�"O8PFN&�bi�����Q���c�"Ot�ZiVd[p�O��E�d"OXI�fO��L���\��41�s"Ot��%E+S�@� ��������"O���W�S�"BСUf��$aq"O������ ���P�\5w�t��C"O0��`늼|�� �pё'�*D�'"O�mK5���G�v賃Ɇ���m�"Op��7�Fj���I(�p�R"O���B�*(R�A�G�Z�I��"O.T�fD�o	���%�DvV��s"O" q�	.0p�Yq���g_(�(G"O���f�P�%J�䉽L�M"O�i���=k9�xv�+E4��T"O���7NP�D�m�$$�/X)H=Y1"O�0yV$���<XU��"E�,a�"Ot`!'���^��0� ��@(p�"OJEx���0A�8�V� �r�B�D"O��	�`ťHǔ$�OV!;f��e"O�jFIшP��!���E����"O8b�Nܭb$��f$�" ��h�"O*)�%oXA�}P���oK���c"OV��clP���Ti@@�0
�����"O�,0�ת��	ht�ûp�)��"Ox5YnG�!����]}Q��"O(�Ⴌ��Ɗ$A�C�3d�P��"O\�`c�2?��!�3[V(�"O��R��:	Ur�",؈`���F"O��k���i8�˚=d|0�"OBUb�O�w�
��#E�t�IR�"Oޝ
vo�ե ��Q4�U�O��y�C�Lf�@��j�I�n}C�& �y�O�S�p� c��	=�f )é��y��s��+q��Ȑ!c!���y�I��]��� l�1��P��yR��N�$P�脒?���"L�yBG��t�n�bd�1$��5�!3�y��v�,y�����h�H��yb��2x�|	%c�f�������y�/S:U b���&^���]����<�y�����Ĳ�ݙ��
W�I1�y�a
��n����73`X:����yRN�-lZd���g+��ī�E��y
� Xģ��]�&� ]�#��|��M��"O5�C��s4��I<nC�, "O2�C��̺3���œ�x�F8�U"O����>-�k�
�&��8"O
�2bG5N?N@����9&"O���S �c����3k�/=��y�V"Oā[�� `�6�ؔS�����"O��I�ϳx����Q�T��PM`"O��`�2 ��y���'�]�r"O0A`f�{���qUF���L�5"O�p6�C�v/t�z��O�Z��l�"O�a� ���|�X����"(�!h�"O�][� N�_L&� #OI&`��"OĄ��ܳ}�pQ�DԮ8�e1d"O�И��&���ቄ�y���9�"O�t$DI(�B�8֨��$1:�"O�+�J�'�HBa��I��Z7"O�1anʘ.�p<����~�:�"O�h��$N�����ET~�.��F"O���� >8쮥8�ԉ�hȹG"Ov��g�֬A�
�c�ޥ5��� "O���R��r"a��j��Y[1"O�a���>�L�"�O�$Nݴ���"O�a*��,���[�x_�X	�"O^|��,���C�еXH�x�"O:�H� #e��u�ԏ
�HCh��"O��yDI-�.�2Tΐ�T%�Ġ3"Of��wj�78�м�熆d ���"Ot�s�f
GQ�0r0Kݻ_|.��q"O|��15FЁ��uwdX�Q"O��t��Z�)��H�=l�ţ"Ovq��.�!(<�5��!n�%�q"O�xQ�iÈp�hef��"�~Qc�*O����L�8�ZJ�+ڛrȜJ�'<${0B8`��h����@�R�'����B�U�;r�au.�z���6�0)Xw�X5�6�(��~��8�� 
䀶�B� Q'�;R�H���<�>�hE�]&o	���8e�a�ȓ)#$"dK���-�gT�.@�ȓ&"�A���z��h۷��q_n��!�D%R�@�����@C,�t��ȓ4b�Q*�Ƃ7"��G���p�ȓ���
g���#�IҦ�м(����vO,I�7��4DT�C�8B����	�Z�Ď���p�Q��7P�F��~l(� �bJ�i�v5Q�L�7�H��b�N,���-R\���r'��|G�d�ȓ��hj4΋�d�%9��.#g`�ȓJ��ٰG�+E�drGLʧm�\�ȓH�����M:A��,j��=3^�P�� �n��S���h��X(%d�b6ȇ�e�(l�l͌�t1�j��	ܸ���I'(Й�l�p��m٧G�!WdN8�ȓP?R�ߌB-3���G���
�'e�����C�!�a���Xt�'h�5��\:���<|eNH�'|:� E�~|��#�1$�9��'Ґؤ����#�
�\�R�'�:��C�ʗ-	� Ǉ^
\����'*���g��-�T�S��M! �&��'|la�� O����pWber��'�r�tl���J4�T$L	T��'��)j�s��9ЄC�mx>�b��� \Yq# B--�t,�FKZ�6�P���"O�s�K��y����XZ�n(P�"O��%g��$��xȂ�%���R�"O��ˀ )�r��VP9	�"O⹐1kJ	T���˒�xH��cC"O���Wgѳ$�Έ3��@��@�"O�*�j�.1�@�ˀD�Q�F ��"O<�_*���ȏ3�@�)%"O<�2J��+����#&]�k$�1�"Oz�#�8q�x����_@,"O��AF�xx��ⅶx �$G���y�N�1;�0 ���x��Y"t��6�yBh��B��4rr���t�A�$��y�V�e�Ƹ�%K�U��%����yr��f�D�X���VG�U��^!�y�LG�|�JՑ��
�N�깢5����y��!���(3`Y3wO�5y��Ɔ�y��05hk�rYD���L :�y��\�����G�&n�ژPg@���y�iSr�\+a�O�c�n�!V���yb@����i�#���=Ə!�y�]��h���Ȓ}�,�E��yG��e�P%�t��<}��y��M�1�y��'U��`���I�X�S����˧	ֵ��Bj�ʑ8QFZ/I�֨�0�'P�� �.
�Re�� ����1��Diy�	E?袁xR"<!�mI�A��ț((xR�Ojr�X��P�5	�)@F�(*��XZ�OT���'2B��Z�i�~�-��{Qn�m8
�1k�d�ȵH�>Y����=q`��>d|h�+Th�%Brbl�f�R��[:�$��U�n�a�韖���H�?~��rqh�u�|\�7j�ȟ��'��,�ҩ}�B">���@3P*>bF0ڳ���N~�I���z����kL�BǓ'�21�"��6E��┌�@�pA
�"p #�;%	�Q��(Q�dܓ@�vT��$�8#��u#B����Q�I 8���'��q+ �'VJ?��?A�4p&�(G/A��t�+ӉPd���hO�>	x�)�ᮡx!���O�h�KM>�y��Y�V2�6�3��O�&���<	s�H�OU��a��C���m�AȩZ��i<��;O��D��B����b�W0A��5Ȓ`|�DP@a����?�(�]a�`�,�.�9�Ń�Z��� �c� ��}�1ƒ�cURE���TV�'!|dB�4"V�4�2�L�<gr��m���� ��'�6��O�˓�?)O��pxkV�۞{�2]���%y
�)t�'˚��4�
�It�0�񡖏4���?4�F�')L����'E�O3:y¤�e�=��L}2h��e�*�ЄuS�Ksk��ē��ΟHi#� �\(
������j�X5i�bŻoP�p���+��O���HĢX6��c��6[��Q�4�T5<x�X#���duTy��hȾ9�R�G~���?�MF���'r�lpn�stbA7N��j�׊qO���O�㟈G����LY6�w�_5�l��cGݸ��͑��
��B� S)l�<���� ��ؕj5��'�f�:-O�����.�~���tJr�.�s$RQ�F�,H�<���@P�1 �x0W�'��a�w�@�BxHUh����R�r�,;�T�X!ѭ��<~���
ق:W`�xo�>i�Sd��L�C�˽B~H4IE����~��e��K�s2៕:]�P��`�K}�`��?)�����'��>M�cN�e"~���CʂA�Pa�u%}��'�r�|Z��L�FJ�5�t��D��i`�JY��
"̘lZX���pNRM�N	���Պ~��:�V�B\����_��M3�����C	�9�$*Ȅ�dI��a��^���`�w�F��߸w���Mn��ItȄ��Tn�\���RS%�%~�<�Є̔#k��-[6j�;\��m>��d!9�8ᓊS�Ek(̋~�f$z(OH���'�J?��O��Ds���&�#B�dDQ�ЗH���מ>��$\
�{֊��_��%��w�c���hI�DQU���d%��O���D"�$�x���f	��9ZH
&�b�"ՅēW>�   @�?�   �  ?  �  #   w-  �:  �H  tV  d  �q  �~  ��  ��    *�  �  V�  ��  ��  6�  z�  ��  p�   �  ��  ��  Z�  ��   L
 � � v /$ �* 92 &< ?C 7J LS �Y a \g �m �p  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf"O�Ya��=!l���Ɔ�b�V��!"O�!)��Y�fx���eE\z0	J�"O>��pg�0Z�2=�C�A�Hy�"Ob\B��;h�`��Ɇ*���S"O�h�T�ÕZ(jܫ� ��+�Ƚa""O�A���I�{"��qReM.v�\�J"O�I��cR�G�Fm+De����(�"Ov�M�{�Ҵ�U���F�T��"O� ��M�g��l�a��8{�Y*7"O�Z��іh��8`�tm�`�"O&ESS��M�,ɠ��b��b$"O,y0GD�!�<�Y#dYF��c"OV�Wc�6�:�3�	�C��:�"O�`y!�������3-�<�"O��!S��3C����ǇZ��\�C"O�V��vA����EE�@�J�yT"OtXa�Ǫ|�t�2&�ۥF<��BC"O�i�w��&dUj��+,1�4�"O���I�tͰ5���߷O�y9p"O��&�(w�̕Z���
P�C�"O1@ŏΞ
f�}KT��}�P�&"O@%����-Zw*�`C�#���"O01#�m�{�0Rda�#�"O� �	�e���Z� TX�؉B'"Ot�[��*Y�~����4[�h�1P"O��@�K�4Xպs-َbF�ģ"O�-��H�l붼�t,�0F(���!"O�����G>�`R+�0Zy�6"O�eXu럋>���i��wf�%�Q�'����r�ܤ��0a��TA�a�%B듳p?a�a��_�����L�)c��j׌�m�'ua���>)�T��'��L��� C)�y�
W*W�����) !�;p��%�HO�0��'x���[J����e�9&&B�	&$n��
aBA*n��Ep��ׅ(C�I{�0���&� nt���U��2B䉮�>I3S��?�F��TaX$3VnB�I�vnqk,��@qt|���U"^�l��$?ѨO�`3�̀#&0z7	R&s�@!*2"O��C�J�;�<�b%�G7~��G"Od��W3
Q&�
W(A�,�j%qc"O��K�+�#7
)$��.K��p�"OM:��_�K����fŇ2��ppA"O��P��5,"E�'���C"O:��D�*Ah:��%�;'���"O�E �GG\%�]#�dF	kF��1"O�����=Q:��Ȕ�%�Ȥ�"OhQ)q�Z����"eHL�7�h�6"O�`!)ƱG��0�G��;rj��"Ori�*^$xi�0�$��"X�08$"Oh�Y��#<h�@�g�1�Fp��"O$�@�U�j��`�杁*�ޙA�"O^|C��/�=�s�
Rg��6"O$i�7eMz�4���8@��"OޜC�� P���0�ԫx#P�K7"O��Z��t�!��C� fH���"Ox�P%�Q=(�:%�2B��{g���a"O��j6��#b�<D�����c����"O4�ŪΎY�� 5�ѮP����""O��B$�1_��U�ְ��"O`�TI	�&�d@H��o��]�T"O|���晳b��Ĩ%G��8Ҏ�X7"OD-�bkԅ4��m٠��'�N��"O�<�6��"A
�Kް1�̃"O�%��\{�b͛����v���"O�T�+ԊL\b=iC䋧.���E"OyI��r�F��UCڟQ%�e U"O��{х�Iͬ���`��
�����"Ov8J$�W�'�Ό���/���"O��{�@R W��%(�h�Q��;�"O�HK�֐8~����0G��U��"O�5��h�<��&Y	k�*�3�"O8�XGk�&q����_�T=�g%D��CĞh}�4"'J�\Zl��`�&D�lpD���<z�$J�)F���(&D��IC�I+�vi��å�� �3�"D�xY�iV'~l�f�B/P�д�J%D��j쟟Ms ����K�P��0D���*iA  V˗��z�d/D�x`R���������*Ĝ�y�0D���#�ɟe$�����!¨�q��9D�lq���(0ְ�h�o�hq�"�5D�8��ǆ��	
aɜ�w5D����aʏ}^�u��Ϟ�u:f�s�3D���� �
��`)���* ���7D�d���Ӛӌ��֪U�\p�.+D�舗��{	T�#b.4pU��.D�� ����=$Ȃ��� ~�R���"Od {CaĸV����HO:!����"Oa��X�O0m��ԕs�ҥe"O�<�U5S$>Œu�ƣ(��L�"O�4��0�`Dɠ�Y4#�fi���'i��'��';��'���'�b�'g�<��#I�e^v�c����M�<�K��'!2�'�b�'�B�'H��'�2�'/���
]�U�iQ��8p�bI��'���'���'�r�'���'���'�X�0dLްJE\�0��(�15�'���'�R�'$��'S��'���'׎<`�
6^"�)"�_�@�-��'9��'���'M��'T��'��'7�m�Wg�"Y�9K�MT�:e��Z��'j��'��'���'O��'oB�'����3b�-����)ˡ�9�b�'�R�'p��'���'>��'V��'�T��^@���P!�F�J�̴L���'"2�'J��'���'�R�'�r�� �$h�q˅I%��:���Z���'J��'�R�'9��'	��'_N�"WbA�&�h-l���ܱKm��'���'*��'�r�'�R�'gB�^�N�.�i$�9��3� v���'�"�'t��'�B�'���'�r	K�G_�`�'(Q�MP�ybbҹp��'�R�'#�'EB�'��'��D<��S�ʩM&n��aG�n��'���'�B�'���'�lPR��'"E��N���6�N i9F\ �˞8����p@�9�O�<�/O�O�Qۇ�YDFF��G�E����&���<���iA������y��'!�\xb!�-p��`�g+]|�J�'��p��A3X=$����x?y0�i��d�;	j�èOq����F <�0)J@I�!۲�'F�dG���ĸ<a̟���ʟBiBr�2O��6�� >?H�v�a1��pd���1O�moz���cc�7"8��#ᔮ^xdc�͟|�I�9H����9TR�-�'E��u�<O��3gH��9N��ȘJ�`�2;O|���D��?��B�i��b�p�Һ�"�'�.���*^8�i���ț'���R�G�8)���5�	�w����m�#䬡�a�J"?��d��~� �)w��ß<�I�LNH���D�j��I�!7@�ܫ��ʐ:�>����OZ�ɾ�M{�Õ%4�҆*c�����?لf��nxb��?o�Z�tÁFjq�¦<a��9�l`����W��<�)O|�N����"�Б*i�!>O�LP���æ��� Jb>��ӫU�KW��:+_�[)�I��[?�Z,����������B�b6�ͬ;����ΦI�����j�Dn�"�r�#���*m��L�iN,�'��$]Fj����O<�D�O�鎼G�4m�TK�-�`��۾n=9�,�<	D�X�%������՟��Ӏ�v����@�۴|cȉ���"58a
���D\��!��4�,}�Ty�9�D-�s�?,�"��S��}��{`5Q�d�ª@-��Rz)��"p�˅#�����dT�?��ͪ�by�Eں� �0QF7B_TY����?����?���?q,O@l9�a�]eN��^/^�:�HC�ߞu�.����Ũ7W��d�ɦ���Yް�/�I쟀n�=_���qg�t�PmcT��!�E!A�H,]��ZAko����}����V�Bu+�<)A-��߹�fk۶'�D���GJڽ��N� e��i��ԟ�����4���3�%%?�Vvź�e��8�R�׿d�V �'��l�$ia��Zɟ�0l򟤘�`��0��/��)���ތ>�Έ��π��L�	�^���PA�Ԧ��5N	�m�����E(,|���� ZF����?�Fm��oԮ�?�5`��~rJÎ �r��=#���]Ɵ�I�\{ī�
j^ ��'kꄂ�+��H��Iy�iA�I�z�'2��y�%�����ѽm�x�2	�����a}2e{�>�nZ0?g�	8�HZh��B(
)��cF��5k�8��x��▢�'0r�fGTy��5�N�d�/����"��#�5<Ɲ+��ײi�U `�OdHPK��RF�d�O���O��İ<5(R�I���� mW� ���ܙϓ�?��kP���'��B�Od�'[�&���襑VX�Zt��[5G��t�.7mݽH&P��#�Ա[��D�OV��bb�0�uwL֪4W�	+B��=��@<"�V=�K�o�ʠ*�ӟ���*�ӟ8�I���I�?ёoFT�Dĳ)|,���M6|^b�)�,ɛ-u<8d��{��'�R��y�P�T ����MQ�:V^�I���� lh#��`ܛV�j��*��O�t9$�Ύ���IU~r�]䟜�F�+3�y�3��.=�l�R�c?�%!�P��@���D�,	����ʓr:���Ox�"�MQ�}{4쒩�,ZdM�O��$�O\���<!��70���Q��?���A������4c�P��'�V9�v�Y����0�'����?1޴,��?m�ݲkͫ'V���ֈY����r����?Sjq2�dD$\Jf��,OjlR�П<	��O��r��L~r]�$���(��'Br�'��}���"��O�R�'��08ܸ��re��L�I��lE=`@�Nܠ(&x��^�XJ޴�?A4�|~�w�@�R #��G�X	�\�媆�SN�`�Fq��aY���]�<��Y*��{�Ba݁�s�%H7ْ��K�x4V<�1�԰U:*Q�'Y�[��'OL��F�'���'�O�(�"�M�:]JR�
S�I�`?��86'V���	�97y-+$�ʓ�?���<�O�%!G��%hn�x�ǥ]�2�
�-�<����M���FM?a�&V������?��'$���; k��x�f�	3�U�	�q!+���$�(� ��- U��<K^=��4O;�r��0y��5��@/T�aƏ$]X�Q���4��՟���|y�˒�4�D8�T�'&*�:@=�s�n�x�n��S�'�66-�O�]����$��O�`mZ�MA)1@���4���k׊yy�J٪}=�	��땉$܌�n�/^[կN��"/P�yA(0� ��� r$H��.A9���@��4���=7��d�O����O:��Ki���nX6f���5�ïV��b�.k�����O&�D!oכVEp>]�	1�Mk�C�<�ϓI����!#* Lp���������M?�q�5F -�i>�3�/��3�O2,S�b	8���\^�j0�@�^�[�����>r�}�O }������')2�'C".��3�ցa�)M>�LPs!-F��'��ɸg^��)�ş�8���h�s�К��Q����X��͘N�r��fI%?!'V�(�	ş����@P�U� �)�B�r�a��� ��-�ud��,c~��� �H �韚L���'
�@"H��j��'*F�E��7y��(3 N �?�AH�c�F0���?�'�?����W��FK^�)���Ssd�z���A��'I��D�Ox�m�����#?9gW�<�	v�pHz���2�v��d��0��I���_�r`�Q=O���҈cʾ��\w!Rp�U]���4 ���D:��E�&��ٛ���O���ɦh������	۟D�4fʅ�Oo0�g��ciPv���u7�@+��ķX��YI�V�����?�i>��	;�M�;z�vm�'�4�[��6F��i��6�F����$8��˟~U�vj���0�p�W���}vD�nÌt�@T�|D^����g���>q��'���a*��
3�e��b���3C�$Bv��D�5F��'+�'j��6<� �Sս2��'Or�[F������h(3�E�/t�J�:��D�B}�`p�@o�	��ɍn����ɬ7W�1��n�N�؁� ��ku��Jw��l�m&�(�͓r��d;���Y�7Ft@{��p�hM���?���[��Ũ�FF���?���?Y���J:��sN�
T��x� bR	�?E��<a���?�v�i�� ����4�=K5j<.��ȢN��;Y~mr�ѱHn	3n�˦��F9!��@�;�y��'�L��aJ�ںo�� ��� �,b h��X��Ȓ�>���'��yх�'p��'^��O�E�%G�4��(�%Ќ*u"�h���i�ɛ_����d����IƟt�s���ڟpqf�L�M�a2�iȖX#�M[��ء���Ѧ��4hJ5�\��Q�c��?	�Sk�8�av萔�N@H�`A>oz�`�f)���pS��S�
�l��D
���ɛ�?a�a1
��ƚ�E?|�fMY�o�Щ��#S�?����?)��?�-Ol�L˯s�D�D,bdj0�� �$�����@����u��zs�������M�ihb� ���2��P�w��|V^|۱��bC&0��ڈ�y�'Þ#���o�>Or���۱�w�P`Ȇ/\�<*H���- ��q�'V�P�B�'���'��tlXM��y��!w�H���y�@]�'`Z�z�$�O �DSN��4�����E�I$ ���	�T..d��Ύ>d��=���Z$y^��XEF��Xf�F<b�oz>�e��ƺ+�Ob`�t�ۣr�h�a��\[��9�0"�ӎ-z�<��9�OX�	�q�Y�"�'�� �,Q4��:�%�;hd��HШ.��'{��.^�d�b���	ğ�S���qg&PP�s�ǖTﲡz�#�L~Bʯ>y��i�6��,�����h�婚O����p�N}"8E`�aW{ e��4�p�)�S�}-0��?����O"�c��>��+�'��u�cP���ɠ���oF}f^UJ��'(�O�b�'��ɣs�4��q�ƞ��A�@G٣{<`�Gq���Iԟ`��4�?��G�S~2�>�շiqb�FfG��Ec^#1l~$Qa�	�H���&<gK�x���*��$�"���_w|��r��� ���M�!��7t_�"��O0p�I�A�x�A���Iǟ��ӧU�|��O.8�TꞖQ^�3f�#P�\�(�A3vvxi��'s��''��D�
��$�'?N6=��h��e\tTjX/'��ɦ�@�4����K��L��.1�r��uש5O���F�j|0���
�4�.䡦8OnY3���?�C��L���ɟĹ�A�ş$��!c�h��?IB(��H���L��џ�������'v<X�e�
�9�r�'�
�� #��9b�Y�Q���8rG�/���_}rme�D�l�ngD�I�u��$�6�֛Ua�H:�MG�Jw<Y�@�'��d	�G܋ {,ahe]4��iD ��!פ�Z`h�(���F��!�z 8��B�������3t��;���&?��	����	�_���揓wV����ݬ{��	u��Y	$b������%�Ms��2����y�Ú	d ��`�8K��9MA�g?h�s�U�xv7MG�@���-{�u�'�\��,⺳6"9>�Tm��'YsS�B�-nx��"O����<Ht�`��?���?��[|�A���d9�bi�Li�١�������1��<!�����|��p|�3.��X`<!��tW`Q�QW�d�ڴp���ʡ�~R"d�ē����ĩ&� ̀��\�{8��r'F�-J��P�.���/\��YQd�O ��`�>��'
�����y��kF��8& r��5�ğ+Uⅺ�'g��'���'�削C�|<i1`�ҟ����
8�~<ɤ�Bq�"`��ߟب�4�?9�E�d~Ҏ�>9��i�6��'5'l�ѱ� 
3%%N�9��y��$��$r�4O���זsP��Yw����R^��;5���$��=�FeZ9i$��--{���#C�i-��D�O��韒����(�9����T�$g҆I��S�7��H��K�O2���ODm�t�'��	�O0lm����Bdo�d�i��!�a�PdY�6z��Bh̶L6�I]�ʌ� �Rצ5��j��ŭ;�q��'�pe�e֫h� V�U�Sd��
�8GK`����u|z�'q��d;R��6�Rß�	ԟB�B� �}8��@>h���F���	My2-]�H���'6R�'���'/��
3�-
����M�6輴S�O�T�'ȸ6�Ҧ�y�Ϳ���M�&P�i6Vx�B�Nȗ6,�u�h7:9�p��P}C
�8v��O�^Q���6�jk`V�X1�B�
k��RjQB$�P!�?Yr�_�1�FY ��?ͧ�?�����֑W�H-�
��Z�(\�q�ӕvm�;O�$^���'�����O&]�'�6MG�T��KK�	a\><�s�T, ��mz�����#�z����?�l��d"���,|1��ק� 2�) ��.�N=@P��;(�B #��'����ƞ$����O|��O ��˄T�ʧKhh��4-ޝ���e���:�0e�	4f���)O����4�|�$���i ����0�V��qC�2����޴)A�,��~""(_�,�O�  3b��,ԙ�i�R���!*�+E,�	�&Ցrt�I�5��Q���'b|(�K�����K�\�Z��?ua_%�ɬ(x�;��@
�D�OH�D�OFʓ-9았����?	��?A��.'=��C�>H(�B���?RBI~2�<9��M�DLy?� � "gP�Sd�<:�5Ƀ���z�d�{cP�` <�~�����|�6�T7�xb��*?����N�<�j���'tb�'��d���ߐl,�O�"�'2�O�;�Z]B�@S]DFl2��;y��oR��y�'R�n���Ć.q�i޵ s�Če��b��J<MZgJJ��`�!��Ř�M�QI�w��<^w���OҐ#���uF���`��J�fT�p
 M�R34��Û>#�'�*%���'���'"�Od<0�.ޚc������8%t��2�DѺ��I(t�PI�`�ӟ��	�D�s�(�'"6�)#�_�L�X���	&��u�O�>��i��7->�������h�ΟD ڵ]
��)"��G*q~�Ȕ�	0"=�x��KL}��VԞaM��G�/�I��?AQ��d���0�#�Z@���ި5,����O`���O��d�<	�%�f�F���i�9QS,Ϭ �`�WnC+{4���^̛��'�,`��O��'(6͆ͦi`TwF��I�M��3c�@{�H�-:�.��,�.W��Y�~\@��i�u��Ԍ1l����{q �'t#z<(c�Ą^C�%kܥ2��\H�4E�'�"�O��9�����w��5M��$�l��`��1on$B�'�2�'�����T�'d~7��O�`�7O�P����M��C�[y^�PS���5E����a� ܻ��z�Z�I�Qa$�]ȟ:��8�l���ɗ�e+ā����l��D��w�h��ތ{f�g�hLкkeK���Ŧ1�	 $���Մ8F1��hq!	���	�� �'�����!ձ0��'+r��yR@�?7�V3���"VΌ ��I���dF}}�{ӊAnګT��	��p��k�>���\�:p`��e���q��e�a�%G�1b�`
�'E��0.��Q���	8X�N��D�.:��Z�Ѧ�p���f�z ����?���|:��?I,O=k� S�>�1�B��ܨ3��B��
� ���'��7��O� 8𝟈Q/O6�[�.��yHs�ʐ�l�pD��~54]lZ$�
 ��BX1Bi�ѯ���+�@�#�NAz���Kl�y�Ӛ?`�Ō޾zt���&�?�f��?I��?����R�����)�0y@�l����V�E�чM�w���Ū+�p�$�O��D����(���<����yw��H��-�u��%N��#k�i�z6�����Ҍ���А��A�����RY���h��I�VN���0o>� ' U�+��̓�-���OX���>��'�!
��'�R��kW��˅.�+9�� S�#0���'���'r�tt��I�����I��%��\���b����l�V\`���!qj(?aV^��+�4͛����~�Iŧ��1륤ۨ7)Bh3a-��6�'k���v O�8�x86/�TB��?�@I��H�2�̅	�P ���MS.� '�O����O8��E��'ܓ�����O@�$�� \�9�$�˒U�V!� �q@�'����'��'��7��Oz�	ǝ�杓<P"�0	b�5��o��&P8�4ЇX� �شg�
����uG��,�Ԅ3'Y�.O@�
e��d�1a�0�	7�#q~�;��/}��O@�XRo�O��D�O>�d���6MC��)d��$-yB���a��@�������?��?���<�'�?tH�6U�����T �M�,��I.�M�i���8�'.� ��N��@A���|���8rP�#K�0l����`Ï�{#.�[�����O�<Ps�>�f�'�<��	@8 ��D@�-�b�"�WJ�?S��!h��'�B�'���'��I�U���c�R�D�V���E=1�L�6�����ٴ�?�GK�|~�j�>�R�i��7MZ�A����́U^�<*0g
�W�P�� �W
i��%�8O���k���[w�ry��S��?~�^k��p	$#�%���a��jӮUj$�'��'�b�O�V֑��w ��W
�+G�&�3���CJn���'���'�2@ꜧ�$�'l47M�O�I:O�CǂۢQήA��O�2�P�C�ޱ������ADM�\�	���\֝˦�A��'�<qaA��*D����E7�fA���$1�b���KX�m�'���d��u�Θ��?q��?� H���+q��8�(���X#�?���$�f��P�Sj�O�D�O���i|J����T�@[(���E$ d�I��/?�P� Yٴ���a���~��ɏ!��[��	:νآL��hy+�m��KdQq�`�g����T�"����Һ�V�Qٟ�Z@�[m~�"�	nĔ3c� P.�YEd*aP��$R�"=�(�`*�O��4�~��O@�p�t��H�O*+B#ɢ ^(��s�Ҧqj��'Db�j���$u��I������N1 dEس�Сy�R��mL?�M3 &��o,�����c�'P����OĺKF$;N����t�2@�ـ$rn�+d��'��O� H��8�-���O �D��<Y�� �|B#(C�}�61�4�0Y��ۅ���,��Ę���?A���?i����O)&j��n�b��0���KH�}��݆9��mZ9�M���h?�����$�BI���?	��ź��4m�6dЀ,C�.��8& �(�A� 4O8�J�!�"�?)�C�����ڟ{B��B�'bȸn e��Z��:b%* �'�2�'�rR�x��͸��T�'�I�E|��A#�<ɂ]h����bMM���$A}b�'��,��~bL�2I z�Y$e��`t�#�V�id~p&jM��?1�LBa2�sA��<�zp��u'*�?�� �˅L]�+oJ�a��T�x;�Q�`��O��d�O�,zR�Յ������d�O���ۏy�)[RK��B�dW �����\�J [��i�R�'l6��O��1期�]�sƤ���Cُj4��1bֵD��E�d�x��:F�����uw S�'vz�3���1�� ��*G#��d�^��mG�n�I���Y�r��?�4ʉ��M�B�'2r�'��$�T&dن��Tw&4�"\ zQ��S�iA뛂X1F���Ο�	�?-���|���c:rH�@$&&*b�E]CT��0S�0�	���"N���{�j��ec�����Z�P�`�,G�l�sc�&r�:�X��׸Lcx�"tɫa��Í]4T���G)��;`Y�,[��O����2�+f��H�)�"rR�}"��������?Q��?����d�9ˆ����O� �K�9f8�l�3Ȉh���#t-�OJ�o�՟�1'
1?�w^����9P�"j�P�����'l�`�h�N�^�`E	eM��K��8�7&�ß�i��j��Β��D�{�'i��I��ru�δu��J'�4[����56*�NIoڱ�?i��?���NTe�M~λtB��{q�$DH��gύ�LIZ/O���O�@�oz>��ɤ�M�2^�-�ډ�����*���r"���~���v�����S(dx��l�O*�	(��t�1s
]��,%z�b@��DZ< �@-����'Ϯ(����-� �'D��$ҍ �6mП���ӟ�Y�'ʑ9����h�O8���A�͟t��MyBA�Oͺ�U�����?KV�`��(�#+�ҹ�/��;
��b�6?��W�l/��Yn��*�Ɇc�2 �4��]�#C�	DN��U%� -^0Z e�13⸨���	P��"G3O�Ԍ���?�hSr�剌tR�L��F�4� 5�G9A����2>"؂DZ�?i��|j���?�-O����c"wJL|�R����K��n�ȟ����M���s���'���#���X����w��&u�F��1�Fo9r���U�n����j������cK�A���00"<�	�'D�D������A�6V�A����� �".C�H�B�'hB�'���
:V���T�B�y ��B�j!:��X���e�䋄�`�I㟤�I�?E���|b�&��wG\�W(*]NJ���[�gK�A�v�'%��ć�~r��L�X�O�`�
�D�̥ Gc�G�d)7���DT9$"�/�y!Y��X�ɗ4#���/Oʝ��)K��l��?a@�F�D'Lܰs �-������ǩ�?����?�����T9v	Q�n�O��d�O��h�nU�}���i&K�v��k`��O�eJ���t �O��D�Ol����O�(���<Zi�Pbvb�0S;ta
�ʣo침2�'t�L25�&!$�����<�yb��X`��'��%�ݍ=	"I�ׇ �Q�'ܙq�|]�IΟ��	�g"L��`G�������͟<q�E���  ��:�v1zd@�П ː�W��MC���?�t�i��G���4�Z�٧h�:zx4Ђ�S��CT��*H �rI�O�x�!��C�V���Z�#.�$O1�k\wl��+�'#��1��YE2!h�� `�'��䞱d΀6�ԟ��	�\�S^��Ū��Uly����͓�%cy퍶zB���t�'���'���y��i�OT@
�KJ�m�  �E]�ǈdB3&^f})x�Ԑm�L�<��.&�\XJe��������FT���Ku�2�����e�L���.��(c<O��z�I�?����50(�I��?	D�P�D�pClE.A̞�7k�v�vT�ԏŲ�?����?����?�+O�5��G�1 ��L+��Tx�"D�'�~)�W��*K��Ǧ���K���+�ɷ�M#��igX���`�.2R��&�Y�IF���է�07&�\�C�n��'y�-p3�캛'�[���ʧH��K�T�E&��a���H�'����i:����O4������+�9�~d� �S�^�M9�~)�P�$h�<��I���ҹ����'!�6��O�h��3OjA�A(An\#W �$F���P�!J��4!�؀-g��ճ*|X#-$!����r�"0�֩�1vdh�i��P:]aLبR���?IǮO�V�剒�?I���?���?���,��v�m�X��$M�Q�B���?!/O&�uL�
���$�O,����2�l�8�0,U�!+ƻ0a��<*#�����$�O`6m� 5���T�n��E�O$̜���jBq��m�,�X����A'8d�T6Z:�xۙ'j뮏��-����A���1*��>�N'ND�q�xI��'k����	�}������'�b_�|��]�6�2�.��-S��;e	Z�/+�]j�ny��u����@& ��������a@��c�t��m0AI�(:w����Mq,� (�n,[6�M3m�� ��:E"tcz��J��3e��tژ��'�+da�ͲQ��B��OX��I~����⟼���?�:%hN�	P�voތ)v.*���z����`�|���%�.���'"�O]H7�<ְ�y���z�	���Z�)R�聵Q�N7m�-�d���n�\���6�%�kv�U��-w�F�ꁤ�;��h�$�1���T�z������CA0e3\� ����)�ܴ1<�i�2.������N��)�k�����'�R�'��ɏ<T@��pő។�	⟈gŐ�	�^ఈ�7?�ZDSٟ(�1H3?Q0X�(��4!�v����~�� �a]B�a'N�|�P� �_yH��I�<�gKI5K�Ւ����f�B��O+k��.�D~�Y`�O�A��Xq��M����D�OP�d�HR���#�+���O����O��r�EL�I[2��@.0P)�vD�O��Y�Φ�'�t7m�OvD�#���+[V|Ͳ�L�7�6 A��ۇ=|�����U�.�Cٴ>"�xuN� Q�+E;����ɝ6�Yw��8�b�?sx�4a%jX$Iu2��/�����'n.�$̇:06]����	�4��3 E[ �����T
�]Y��вo�ryr��f�t`���'�"�'.���g�P�Ix��� �B�o�N�2��Jk�0JW��3�4#B��	M��~��H$P�,=��'���b��_۸��N�|��2�
�Yb���=&ǒ�ɑvO<����'\,5H�D�<	�'����geB> �X�q�M��I�n|:v-��:B
l���'���'�b�'�剢�T��g�N՟�Ƀ`E�"�����G\�,��x˵�a�cڴ�?��j~���>��i~t7���i��\ɡ$��v�* �E�D/Ɓ0�s?B�2gM*n�����/��L�Yw�~ab�@�<]w���A���%����Hl��C�>�0�G}���	Ɵ��	�?�*t�sމC�%�M��.4o�HlR�`xy��'������e����O��mZ������u�p2P��7=JpI3�O(G]����i&�Z�	�Ƽ	 ��O��01V����j�-}5�ē�R$� �m0�&�~HX1ʀ͍�j<���`K���?�G�U�+�I��?���A�M[��'���'�� ����-4�1r.���f��A�'��P��jP�)/)����ß����?��ڴ��H�Dɰ+����M�r�4]�'�ꓲ?i��O����l��pU�Pß�ZiT-s�&�h�h�=a����!�<^�Fѣ� F�4��%x���;.���	"�>m�-OF=X$J΢9g��ؠ�ŠL������SƟ�-D�W*}X�$�O�I�OJ�d�<�Q��@���!�>]���Pe�ij��i��',6m�OP��A����O���W%&�m����+O�̔��3�6�dٶ��Q�NT�\�($��OU��k���u�G�/ Z̰̓'�"���S��4dc���5e�=�	��?�5г�Mc��'tb�'"��	P�Ӌ2��DZG�5�W�üU� x��Ó 30N��������?b��|z����w�٫��ݠ(4��V��#�tw�'�"@��~r�E�Q+fe!���1n�F:И��X�{��	֏�9x�hx���v�ϓa��`(�+�O~����ZKyr��Ol�2�#bӚ��I#d�n��IA�+���A�+�;`����ڟ���ݟ@�'ZD�gm�"u"�'�b"��9�T���Ã&%�Di�a�6*BH'����~}B�'�� �~Bb�$8I[��m]� �,���D >}e���?�1�X�D�I�Q�Җ{R����u�� �?�����vP�A���E� u�V퐒x�F	[���O����O�����P�~�䒟�d�Ot�$����q�gHR�\��Y �;���(XS,�l��������M+��R��i�y�k	&FI�E�b�;j=ܽC`��i�NHBB:8mL7���J�N�LYh�����O`�X��1�u��ё�x�C��������S��l3���pyr��OHUH3�d�Fy��ڟL�I�?(���L����W!ؕu���Z��'f��b���@����|��/�M�'�?�.��H�`�=^�|�l�6i����p�ɾ9F��I2ٮI"�?�:"+ϐ,���s!H/�CB�@� ��P����r6&�1+T��B�'�F<{d�<!��'B�rr/�>XJ�%b��x[��dCZ9yР�P�'��'{r�'o�I)��BD�W�����%$N
^x)6�@3=�♠UP۟��4�?�gaa~�>���?Ic�>���,�s��m
����
P���BH2R�P�EJ�#�?�rm��ם*Ѿ�3O�����; A�B!&oT�G�6���LV'l-��E�i����O��D�D�eF$�9�:��q�%��1g�*L���@��O���O���vE������\��4�?���<itb�>s0�U��l�^q0̸�f��D'^$��ʔ�v����$��R2 x��V�����ɣr;���B�R�>���u.^>��H�m��,��O��T�,�r;�$M?�f��O����O�Z�+�/,j��9��\�m�"�pcf�O���<�!D�|�� ����?I����W�i)�p[�ܟ|p�q� �ie�t��ON��'��'�ȥ�'Ԯ�V�5�?if�׎VŊ憛&Ld��b���E~���
��eo�I	c���<A\w�Ĺ��nO��jP[��󣌪Ib4d���H�B@��ǯ���?�O	�x�V)i��?�'�?����dH P���s@��=g�����I&|i�	�3������՟l��4�?��	�]~$�>���d9%���$T+�*\��$���H"�S�.�,?�@�Bw�\=�?	�G1�.�'��%��7Od�ȲL��Jk�P9w�#-bys�'46���J7�U�����\�S"����O�h[u&�Xh|�i���^/P����G�uѠ�'�2�'��T�zӐ�d�OP�4�z�bd,[
:�`̛�(\C\�?���̓yup�`� ��?q�'O
� l� �Ƥy�mE0��ykb�\Y�@Lj���<��T,G��D�	V�p��'޲����S�Z7-���<`������f׬8�pD(U�ҟ��I�x��Uyb�7E�n����'Ub�'h8! �%"��U�2+]�	P�'���O�'R�'�N���'�qQɄ.z���&@z���h�9����]�pm���ZQ�BĹ��D�<�]wd�9����,���=.�|���S~�9�
�)�0�$�OP��$$�,�˴(>�I�O��4�hc��*��c�"0�|�ug�O4U�7�����	x�޴�?A&����9�Ƭ�����/��U >d�$�Rf'=Ub���)ʷ���b��Ps��)S(��#M�:UA��kl��`����l(Z�9pd<����<Y7�'�����i��D�O��⟔��bO�5���r�"^�x�;�G��(��_�T��8�6ؖ'���On�6=���$�\[�yF-lE��4f��$:��'h7����g!�� Z �D�{���6N,\��m�Ĳ �u�5�H�U#�>ܘ�@��e��1`�^1�ćL�X�R^bN@cH@�;ؘR*��U��7@��H)��Ȯ/�R�'q��'HBY� �7hև|�\0��8o&J�C��@�=���C�b̖��	��M��#��I��|Bd_� �	��F�w�Dh���H�NX2F��rX���N2`�Np�g��ퟔ�b"��w��.X/���' �����9Hg�*D���  I �( �qj�) ��n��?����?��'G=
�3I~�;$��=Yg��!T��bk��0�Z��?��7�̴K0�iH��2�M[��0�"�ϓD�x�s��k�z)@��!ZE��zq��X?	sG�il�� ��|�7���{�z}� ��<Y@ϷN=��cFA�^�i�U�6,(ѕ��OJ!{��E[yR��O�t�E�y�Z��	ޟX��$r��	�A�( �&�ƊҮ�X��ʟЖ'�:X�	~)R�'>��O��6mF?O��-	�߲*��1gG]>����D�ܦ���4tH��W�aۥ�f>ex�l�3HH�FO�9?�F	a2���d��c �h��ER&�v����!>8B�7=B\˓Y۴���ȅ��J���q�d�;��Ɨ�\�� ��'Y�O{"�'��:r,�Ō��8a� �2]�1��G �M)O>�n�@�-?!�[�(PܴS���@� �7fo� K�"u��쏜C���"A�_�Və�@Z/S��;�',����nѺ�&+.7��I�"���B������ T�d�(�����ɦ�����?a��bp�Ӏ��yfqpG�[�K�d3`��h����:$~����O�����o�wy�E`����p*x��g�� �@
���T�4m��M���a?a�mA:1���'U?��`�!��\.�� ��@��6+~Iᰨ�#S��� �8Ol�#S���?IE�Tpx�
�?�$�Z,�M�U�'��]s�bZ)I��mB�A�A!Pq2��'	��'9BS��hǍ
�R�2�'��M�r�\�7A	���	D� ��
� ���HJ}�NnӦ@lZ8�6���PHE%�/$�ڕp�A�',r����-
���d�$S���pEˈ;��HJ�^>�cG��O�(��;@�z9z3��6TwbT�Q��t����?������(#D ���'�?���?92�
=d|̝`�}K��ܞ�?�'$_dꛆ_�p�ڴ�?)%-�C~�w�v�gػȨ�a���C��qY��V�7����zӾ��@u��2��=&���V
~A�Zw�$��e�W�^a�(xW�M:��A�T�
0XK~��'���D��
b7M��|��͟��=�V�0��R�Ox��@�_�:G��k�� Ay�e��|(�_���I�?�*��|z��<��P:"���3ѭ֮H��y�UX�8�	��Iڤ(�����ǒOV�><�P�Q�aP04"X]�D�\�5B��ˉU�a��F`�`�f�N�D/��J4Bn��D��H��aaL`k��)Lf�<i��?@�6I⡢o���'Sr�'��'��\a|�2 C�؟@!ul�	S�A��
.���Fԟ�{�4�?���[~�´>���?�BJǱU�,��r��3Bo�A��h!��L-�>  �
j�(Q��JL��jb�0�B�m��+տ��.H�{����'oy��ɓ��R�bɱ�46���'2b�O}��W���w�f��Fu_�؄�C�_��:��'f2�'PD4���n����OIoZ֟3�fp�,��`�"��9!���l1�m�fN̳[�>�I�/S+@���O�ԬBu��?-����'ɖmYf���r�� ՙ	��	 d��Dq�|�I�F
z��)O���	<c�,l�?����?��kܮ�p��n�&�%����?����D��Gr��#ū<����Ųin�H8�jܸT�lU��A/G�d�h�'���>�2�i��6m8LC���0�� I�OT����O�4 r�!n�����#��?z�L��=!3d�#���ŋ����G<���d������9uD�� �	w? 0�I�7���Z�j�|�i>�����,�'q�9!�욕j�����jź�VfY�{ʼ7�O��D����I�5fD�d��I˟؊F�D�u�h�i�5Dؚ=��%�ş[��]�F��4$oއpK���0j��9ƹ��CO��y��Z�IA=�r�ŋ	;��������?as�'F�%���i���O���� �+�|rg�t��.�+�䘲 ��oh@�X�j^=�?����?i��7��Ο�%nz��P7eC�h/ ��
;K�q�@̤�Mk�iƺ���' �Tz�ǉ�D���u02����]��(����]��!��6�. y�'�p*f��<�$���D�ٟ������9���'*{��ʩ0��i��J�-�9����?����?*O�����%5�$�O���O�^J���f�U�gaL�x���ȶU��	.��$�O�6Mg��DD�S7"qCi� ��u��N�W���*rf��y�Mͣ;�Tz�i�F/hp+,��9O ���1��5��-dq�0�BV=�ʑ������I',���N]�����	۟���0��4��ʺh�RIŁ���l�R�\2�M{/OJ�o�ןDi�h#?�;�� ��ʞ� ѻc�wB��C@�U�'�r)IU�itNa�gnȬR&�e��A��y��}�����ò$��fZ0C�	#��rd�ԃ:X��,O؝�I�Q��l��?q��?��'��0�%āVS���5��Z~@p��gT���P;I���rҨ�O��$�On�	�ٕ'����ҥҫel��2�i��0l0�Z»>a��i�7�ͦT�$n[����O[����@L���|�r}sP�ϻ\o��B/��μ��'3<�;�ĘL!b,���ӟ���]X���N��d�$W��9� ןh�	��	ן�'�V�{5,X�x^�a\�l�8S�S�R�FhYR��7�g�F��ڗ}���"����O��d�6�� b�� CV@�"�	߮2�̕�de���*�4,w܂�$Z�eV�(Zw�$qQH�<�^w����O3	����c!�*�f�	��[W� �K®~�l��	�(�	�?���B�s�=��ի_>�U���S5-��0�GYӟ��I���#3G��M�O~7��O0=3�2O��3��1����ӎ�&����[���V?6p\u�������!d�j����y���f��Y$�	�l��Q(@!ī4.�BP��ޟH�J���^���jB�[�a1���?����|�`�'��(�p�&Co�����?(O�qcI����O�����mZ-FRJ���;�J���ƀ>P��r�ߟ8n
`o<�ɡrU���1�0� ��f�l1��,��H2���
D�&�0��P�C�Y3;O����?��aȄ5��I< ��0sk��:�Ԁ��l��YH�%^p9��eL��?��S�I����'	|����p�2��<|�|I2 ��7��O$�����	%d�"�J��	-�M��n�-RZa3�m�|�����_�x#
+:�X����O/Ɖ�'>��S&�����V�p���ɶ5*t8�aмFl�e�e���./`�D]Ɵ�;�֦�a���?Y���R`*I	��)@����T$/�2�`�W.B`��3��0GN��?1�'zǛ�O2�i��M�x��!�%% ��H�C>3P�oډ�M[5 LP?��ˑ|D��S�?��b��|�]�R�Q"MZݱ�&�+&�8k���]�(�IScn!BZa�M�l�4�$���4*/����O.��ql��"װL@���-�.�����O��d�O��D�<��w\������?����SdK5%%��W�-�5�T�J��'�Hʓ�?9�4Zs�A�g�X����2]dY;�R#j�}
���b�J�	49�"�;'��* Π%��|z3l���C�wzV=�I�Pb]���¤I��d���'�B�'7���f�?G�O
�'{�5gj
D"��ˬ1"��g��2e��K��6��O��d�m��U���ӼkҶ9���R����Y|����D�t��h��4��2��ȋ-p 9���E�<��k*���]�J1x�"3,G��0tA��&L�ʁ�s��2��	��?�$m��M;��'$��'��$KַjFlS���Rׄ[@�0���
��$�)�$�	J�O��$�O��i�ަ��'���%	F�n����&�2U���AG�>�Ծi�7����DI*J�U�ɟ���!� l�:������c�k�dr$@(�LA�46O���Ƃ��?9��&NZ剤�?�(%pf�� 0��%e������Ѻ$G��8�Z4�?����?���?	*O�kS�m����\�Y�Pa3�9_�ZL[5$3fF���O��i�	T���R��	�MK�i���it�E=}��A
Q%�+�r1�a�4I.8�w�ƿx ���'Li0��������Qp �	Һ�F�w�zM;�+4k�&��e�W�,_��z��	A��f��Ov�D�OJ�i�6osx����\*���tJ�%�V(��R�'���d�O^��m(mz>I�I��M���<P̓q��p{�k��4ꞔ01OV�~��	��{?�D��!�`A��4����!(��Ssi��?97$7w�8��G��c[����&�40�ר�O�Xr�'�oy��O��e�q�~t�	ߟD�	�|Òim�<#^��+�c[-Kqrd��Ο��'�P��E���{?�I����ӽ�M{��H�;�:	3v�þ�4`ct�K~���>af�iO>7��"R�䔄�@����O.�y�4��$��B�%�@ �E�#J;J��QoR�N#���'�n	��d��N�J����#��M���A���.�أ�'X�P��K�E�R�����'�r_�h���R�C�ݢgʯ��0BU�'-���sܴ�?��/����'�<(:�O
��'�m�)]���j�KF�.<F�pIE�!�B7-�`]���?h���0�O�m���Ԍ�u�Z�o^��ϓHQ����	�1q��(��J�< �	�	��?S�	��Mː�'�2�'�����6o�S�P?���AeR9i6agJ�M>���f@*+J������	�?����|�]���wj2lSaE͆� �a��8�,}���O�6�SD����Q���ؑ�O���'�".�.}apI�"R��� �GJ"�:E�礃3T�Z���'*l�6�S�<�Gl�	��D����"jU��	*P0 	zTDݢ(i�Q(WB6A �����p�I͟<�'�b��5�׮1��'�OI�Պ�TZt���h���=Q��H����O}�h�
Eo%~�P�	$9,`	���μgܮL[D�)^����
�]��D
�,P@�*�@�@8�7_>�P�q��I��$x��7@R�t186�K�c��q ��?��,�������䧗?9��?	�,�L�X��S���� P�Kݜ�?	�;\�6S�h�4�?9�,�z~�wsJT�����������/Q�^�3ǘ���W81ԛv�N=yJ�Y�ӄD�>��`�'N<���j���+�� �n鑄�Z129�# �[���`Ȧ<1��')4QA�i���D�OV�$��8p7 U
{R��s��soZY{��Gl,�Y��¢�τ�?����?���-���T���X�a^�h;d��rt�Y�o�7��Dk�zD�|���yC�Od�J"a�����O��S(w���B��<{�5�`���o��B � .�yҧR�w�bm�	����by��Ok��}J�iy��Y#d��I�w��<(V���l�2�?����?����?i(O��(@	�f�����h��Y��Ρ1V ����U�s��Ӧ���7y���E����Ms�i,.���
;fH��0�KE8���(ڪUKS@�$�DUP���<���5eP�ם�V�~\H�R>�h��;X�������b�,� ���H�����3�?)���?����%�*��缻q��B3�E��B�aY����4�?9���?�wfÛ�O���d����Ɖ��$@�Y�>Y��� �V8��+̓�`��O�i;�Âv	6=�N@au!ƻ ,@�cs=O@�u/L�+����wiߥxpƜ�(�!W�4����l���\����*��L��4wBb�'cB,ӌ�@\��Ǿd�N-�§F�2�'q�	02�L� ���������%�M��j���I�gB�)vް�lDV~"��>��i�^7M�)~����6E܄��O��m�k�u���$�I�Ld2,[�.ȴ����$�K^������
����������|وT�#((���)VB1;�l����(ъ��.۟��i>����H�'#��:��fg�,���u���"'K�||h6��<q�i���Ǒ���s}��gӾݱ&H�v���cw��f�Uq �Wݦa:���M�8�*�%"o��'/���W��H� ��C?y4#1�� #�KT�)�"�)5l��
��mڀ�ڴm�2�'@��Os����[>!��#����D'G5�۠�\.%�<��؟������3�M#+O0Hlz�{�ß,�ѣ,�
p@�fU��M���ik���'(,�S�f���H�8��c��%k
��q��.�!1B��d�d�0�'8��7�PП�@�	�����8�AhY�͓L��i�6�H�lډxSDؿP����ɻ~���0�[yR�'q�q²ܦ=��
2a�3�'���9�O��'M�6�K��5��̢�xئ�\�5����6������6|�n�a?O�!s�S9'Ji�'�Ӱ5>�S]�^�鿃�H����£S"�A�U%x�61�P�5�T��`�Z��K��D��u���ܟ�J`J�r��O���Ǧ���-,C�Ӽ���4�~P����W�x%����k���Ф��j;#����uS����'���0bFCԺ��[���r"4LR�Y��-f�8�{!!ˏ���ן<��Ħ�<ͧ	Ӹ!���T�Q"%A�������QN~R����<))7\�����?%��t��m��~�+���sT���uąg��A�Foy�ʍQ�O��� �N���I!g�Ls��G'X�����6L�T)����� ]�p:E4O���G�#�?q�$ĺS4剠�?�A�ÖR`�1g�ƄsI��1�Y�i�N+�n�u��h�ƅ�`����I�Y��UI׊��,�%�e F�Q�H��� �M���E,���'X��%-��At����0� �s����dY�'j��-R@�@5#��}�6�r01O*�@(��u�Ο ��O�nC�'���"A�p��A��ř�)�4���lӚb�擙S�F#<qG�ǩY�61`�K�+X��1I1@��?����?1dk��
�t�t�v��$�6\h�DT�DR
�q�,�Ǻl�ѭ�gM@�8��On�� '@�@�$7=�HX��	�DP3b:OL�"�*dZ���q��&Hg>��ץR��v�
�~����]����.���ڴ^9b�'�-�3���װu"�*��E���'T�ɧC�P�v.ϟH�	����� �M��ѦM��ęV(�c.i���b~���>iǲi�:6m&-A��W>�(��π �@��F��bT�"޹?Sv�1P��(���A�k�w�~��c:O�$��?�G�O�?��I/.��I4�&|t��r�Z?}�L����w_B]��n�5�?���|b��?Y*O�H���^�.'���,�!-&��!��v��1nsyB�~�~��ԈJ�ɇ���Ȧ�ذ�B�N��d�:���W�K�M���܏���bV�n=�{����cI}ݽ�4�V���قp��Ѡ���)eQ��
�#	�Q�"E�OHl�bFxӺ���������?�S���[��֫;�jвb̈́�n��PҢ�5_�Uh2̶Z���'v"�O��6ͺ<	e��yw`ͥvj��Yr��t�,� ����O��6M��xϢ�|�ŭ��I��S�5�Z��&��[�B��yԐ)B�����A���U�2n��	�{�����'g$�+ব<9��'��q�il��"E�"��m�J)Xg�Şz{����O���O�"��A�E �?Q���?)�GD,6����
��-"l|�6H�$�?IuF�}~2@�>IQ�i�P7-K�)W�Kf���H�c� �f��;N�aI%�-�yR��a
��0�ݕ�(�P*�z�h��'X����9{0<�bc /Qm�դ	�d~&=������	5P�T����s���������[��EB���B�0,d��R�KT����5낻�M.OdlZΟ���.?�;c��+b���$�p���R�'�t2o0�Z��a�i��-)��Ʈ_��mk��y2��bl4 �;vԘ݃2�[e0LZ�K�Ou��q.���n�Q%2��Z��v��OR�$�O����� A�)z�<��Ȉf\���<��ѧ5��X���?!��R��i3�Ih�\�$ eT� ї"�!k�zX��OX-o��M+TMTW?Ig�@�R��'v��4�	�����[����Q�mSj҂"���<I�GN�&�$��Is���'f��D*|��p�&�i
NŒqJǜNK�|s��M�����O>�d�O����<q�U;{;�( ��l#�	ԫL�:P�.�D٠�K��)��6�';�|c�Oq�'[�6����x@J�{��%R@�`ye��ϗL�)
FD\�2Nd�*�t�d�T ��y��L�L��Y,�^���7Uђ!�G��4C�B�&"<r����C�� ���?����7c���缓F��-^KP}{6�Fma�ECP)��D�O�}	�*������ٴ�?�凁�<��
N�$1�y[oR{��<�p�YN��-�y�~y�����M�'c��o)q��MGpŹ���I��=�w��<%��W[�����c�p��S��H��3��)��4}��'����Pz �˳Qׇ�,ZY�	՟��'�� Cr�˃MW�Iן���)�M���]s�ѻSJD�H3,��A#��<i��]��͟(l�8�<��4p�B=���Ҭ���I��M���֞	��4�G{�I�FK�(�Zm3`5Or�]!i(\!K���K��q�)�+�X���Q��`�W�H�1F�C��P��L�nɶ!AmHt选�}�l K��|l|�p��H/���85*�8�����@/��p٢n�]�'}�R���
k��
9Ffl�Ҵŉ�H=j�`��8����FS,I��j Ү|&�i�B��u}� �Ō�r��Z%)�\��7�ӥ����@X%U� ��c�^��c��,��Aq�F�n݁�LO5|���)�}��j&�p��b�<�0 ��'� �
%��N�UkV�ߤ�~(��iH���/.�d�O����O�$�'
��](�NA����?u[ ��C�:�^L���'Q�	��D���@�'Xl�e>� ˚�!tbD�菗O���C�y�nE�>O��V�01��Ou��'�r$2b�O�� �	�ӎ2��+;���q[���	ݟd��Ly�$�9 ���'�?	��Qd��@�̜!�|I ��4����'K�-��'��d��?�&LL��Faq��N?%$b-(C`>�\n�䟜�	ly�#ڏEK��'�?1���E�4G�P��a��u����;k���x�����ȟ$��b��l'�Tk�wɰm&f�n�4�8��W�M�]��4��DN3-&x`n��x�I�@����d[�G�u�2��8X��$��|fH%*���O��d̨fT��`Ei/�$_gklp��J�j��1K��ɹ`�����f�P7��O���O����j}��E/�y�oM֎Q��ΐ�b�*�5��S��7-U?2���T�6�쟬�&�$\��daQe-|�)���^��M����?��e��ES�`9�Oj����$�(\9L4�6M�f�T�)�X�r���r���?���?a���O:m�׉	-:�
]S�=g����'MV�{qU�,ۥb0�ɝ01 ��k�� "���/�'p�'�_8��I~�0�$����֟��	~y�	�@	�ij��������I=S+�ȡ�R�����柨���/���6�d�O�x����%P�ș�5D�;,+*%��j��z61OJ���O����<���qP�-_�"9r��;s� a�p��Y(���΄�yr�'6TH��z��?����~�oӕ+A�K0c	/g�0�a�������O���O6˓GK�u��\?}���+�Rh�Bd�N��� ��R��Aش�?�B�Y?�7˝ޟh��d&���=!G@�*��� �R�y���`��K֦]����T�'{<ق�b�~����?q�'q@�Q@ D�S��xI���cԺL��K?`�ڟ�I�k�0,�?��3 v� ��Yh�(�%����бi��8oW��#ݴ��Ɵ�����]�����M�<�!��Q����CP��Ԏ�ȟX�)�S��4yN��1c_�2cze��	Z���oZ�}���0޴�?����?9�'i��	�BM��\�d��!G�֊pܸ|KB�V�T���l�>c� l�Iܟ�&���<���T�\� �%�
dh���׺$l�2��i�R�'�Ȅ<�˓ -��S�4�wIiӾ)����*k�p��BG�Z6E�i�r�|��~Γ�?����?���~G �Ҵ��
_%����@�0+V���'̶ JaŤ<I`s>1�I�S����,���^"O�d��a��;�Pzf�x��'�'��s�8�	�ta<���+�&>#�1C����P0��Ȝoyb��6^��4O��~�'�?a�O��X�!aF$�����?z3���ٴ4��1�<������O����?� 8��)Z����D�O:̬���i9t�۶�'B����~�'�?*���i��St���;Ԗ����Q
���O�$�O��Ľ<Q�G�W�O��J�Њ�l�u
��4����f�`�� l�dI���i>%�I��''��{S��gᄴ�X{d�����i�'C�	= ���:N|2�����sKz��w
�Lx	㈒6��Xt�O8l��[��Yw����9O뮂�-��s2�M=�b�c�LϗD:��ӟ<�5������IПl���?	�'[@���N�#yR5Y��&#B��35J��.O�7O@RѫG��O�O�(�d�H�n�
�ښ^3d@Q�4xV�����?����?�����dM1n��i��'\�å���3�F�R#�]��6��	�wR$t´�)�Ɵ�`������ �
%P�رk��Mc��?��aM
��wQ�Q�<���_�`�v��a.l��`F >X^��珨�M{����Ga�3?��~� ̧l#��r&`��8���
���Mk��dO [+OԱ�d:��I$���O����g,*B~��+G'.�Rt@!�ĉ11�����p������'f �D �	6l"	�"ϔ�y�4[�d��3���}��Γ�?y�
@�<����?q��Bъ�k�`[[F�lj �Q�iG�=#���<�-O��d�O��D�<a�.�=F��w��� �4���(��7E�f�±�y��'v�p'����'	�ɚ�5��2�KwKǲC���1���Mk���?����?�-OR4a7ha�$��5�b�\�����.$r�x1�LY��M���Smt�̓/�X!A���?��^~��Mke���#�"�$O��ő7$�̦��	ʟ��'#&!�po�~Z��?Y����b�f�r(P���K�9W��ȃ��<)d�?���mr�'Y剞�y�`/�)��ESr�F���$��M�*O@E���Φ��Iן,�	�?5ʩO�,��B;i����⍗!UH�0��Mq(�d�O�3�6O��Ģ<a��Y�ӝh�$Y��b�D2�O�e��7MC�	�o៨�I������$	]�Ě�mE���Td�9q)�]��l�[}to���T���߀l1���Ԁ^��#4炔2�<P*�̻l��5lܟ|��ǟ0�ƣT���$B���O��Ӻi	�D	�L0����T8#���ڴ�?q)O��s�3O�SƟ��Iޟ@	W�CH�L�@!�2��ɹ��\��M���g*CtV���r"y����&v��	�?ט7�䍙��.�(�$�V�^���)!�=͓�?I��?Y��?�.O�\���:zQ�X9$͉5	� D����ȭ�'F�p[�'NrO�#�yr�O��'���	Ĕi�lj��V�4	bU{��F�y��'��'���'��,zE��Oʞ�¬@�J���*�#�zc����4��(��?ـ#��<)�'�?i��̓Af�db/>F֍�0�E1m�LA�$�i�R�'IR�'��I����4��	R�:,�u��K�����fZ15Z�lߟ��Kq�H��ߟ��	$d��vy`��_9�@��aߦvA�=� c�U9�6��ON��<�cBŬhl�ҟ��	�?�x��(i��CW�ٰmS��W�C;
?���?������3׫w���	py�.iީD��<?ڑ�1HڂE�q�C�cӊ˓N��Y���i���'��On��b8&�P���j5h� �XHAs���?���en>0Γ�?I-OF������60u:��YE��hE/�:�M;���0)��f�'.��'���J�>1�d��<FĻw4�q����0��)h�鐪3�fŌ1�y��|��
'�O�
�x��1�d�ʞ�^��!�`�7M�O����ON�!0q}b�@��yb�'���B�4���Gd�X�J�G�(Sr!�>qa�R��?���?�w�̸n
D���t�PT����.'���'�$� ��>)&�<���#�e���1o�X!e�#Yȼ���a�<"5�l�'Y��Z�y��'vR�'��ə*�.Mzg�@�p�h}h�,vо�f#����B��D�O��z�1O*���OF���*~PE# @��1�.y2�㞶jЦ4[T���O��d�OF˓��q��<�N�Y�JQ�)5�� �Ȁ�d��M���ic¤ �'%�팸�y"�ORB�'�@�'`V����Y�%#�L�j�V̠v��>��?y���dˀ'JD�O>�ŕ�+�f�C��_�s=�Ւ�[+&t7��O~�S�2O��� ��OJ����ϓ�?)�'<1y�b��|Cʥ�-�$QUj�zݴ�?����d\U�H��O�2�'����]�1����c'�/T����Ӣ!�(T��'whM���'��c-�yR�'��ɶ�y���2Z�R!S�B"/B�	�i&�M[.O�)1�n�Ȧ����jӠ�iDH}�L"kɂ�[r'��mʼ5���>�81��'vR,��y������'Ʉ�O|��J܀' 9@�jՇ3`���/�̦!x�	��M���?���B�P���`t�Ί����00�p�ACB��d����iH^p��OJʓn���|J�F���cf��+����SZ���2��ij��'t�D��{�2�+�ʈ��?iW�ئ����g�`�I�
')T\<!��{Ӽ�O`�77O�S����	֟d)f�Ң6���4�p^�aô�X�MS�0�x6^�4��Az���44���	�?�X o������*ɒ)��hQ�Qo��R0L͓�?q��?����?Q,O"�+e&
/QZ`)���vz�Re��-*R��'ݘ�8���?���T�d�'H� ��)����M0��"��L�*�����'��������̟d�'A��TEn>=�BU�s���K�`�k)����ÓI��'o�CJ!�~�'�?q���n���0(�*��K���E�4s�	7^�H�������xyҬP�vp��Ȭr%�"�4�Bv��X鄄�7��a�ɢX2�	H��$�O�����O��' ���ڃ&�2Ej�˅r��	ݴ�?����.F9�A%>-���?��
� 0 � �B7k�����h�	�nL��hB?�r�EԟL�ɢB��U��t�ɵ�y��o*����n|��VM��Mk.O�!R����񙭟 �$��q�'d�x�����C�rA9
��T�|��Q)�(�?1�O?�xGxb�?��>S��J��٥Z���ro�-���oZ[ʸ���4�?���?��'D��I�A��$�-|���+I�<#�.��K�%aø�nZ:�p�	d�I��b>e����Y����Њ��4IЄ�R��fӦ�D�O��;)��ؔ'�|E��?�#�V��#݁3O�2s�L �	=�M�I>q�mH�<�O���'�#�(���Ӄ	�9��RO�B2z7��O�9�!XSy�琙�?�hc�]��5&��G>ttI��@-6�apa�����dĉiLh�d�<9���?A���� d��(��ޯCd�`��{�<�Aǩ<y�b���IF`��'�?��uİ��6m<���@�d��?� �s�$���?�+O��$�O��<	�FD6CI���.F
Ҡ��B.�:7�OoD��?)��{����?�	���'��w?���1�j�0����~*��;�nFK}2�'���'2剝O9���O|�A,=j�(x ��J��Z��?Q��V�'��R�'����?�� E4�?yK����O���v�;tq�pz2�|�����Ol˓��������'���N����|8nC]ը=��,p��9�'΋������A����Iy�ɲ�yWFC�
bn}kq钾k�n��6�M�)O�#u'^ئ�c��������'Y�h*�aZ>F�6��BM�!'��¬G+�?i��y���`����))�e%>���F&(#�"@	��Y6��tӌ�Rtf�¦}��͟����?�I(O����'`���dI�d�(�
���i�����v����C�O��O�pW���O*pK4$TL�P �Z<!�P��A���5�	ڟP��'��*,OH�ښ'�R�ӹ�Mk⮀%�zdZ���-n�e΄�$����	�ħ�?)���?!�������0'��$��������t����'6>3�'B�˅�~�'󸬡��Ǣ7��P���*�n�[F�xR�؊��d�O����OJʓ`^:�-\�vm�p��E��MC�cC�T(�V��0+�ON��e߆�g~�^�V^Բ�W7^�\� ��ϔ�)�y��'�r�'���'-��1��'W^��c,�zD�������Pv�eӄ�)�O>��S�:��O@�9O��AZ&�M+�FF���*�i�J���XC�]R}b�'�'��'�Д1�R>��d�,�d�τ!�ԩ0ל��YmZȟ��B��*G#�O@��N)Rǝx�ᖮ>��@�4y,��v�6��O��$�<	���1)~�O���O��H�b
�p�`z��ɮ���ܐ+5�5;�'ٰ��'}ԙ�a��J��c� �*5"�hQL�R�ҥ�Y�	��i&�_ß$��ğX���?}�	\XS� �[�X`S�ըDY����`�����<���C 0#<%>9���W5�(���3������kӆq9�.�妵�I�����?Ţ,O��a��'Z~� JA�a���ۑl(?��Q� �{ӆL���	(pS�c�@�	!pm�=��d��>n%��쎓)v��MC���?Q��L�fH�'R�Tٗ�O���
M�6eܭ]�0S��S���P�a�����'���Џy��'��'�v�C'�r���� �m�����v�b���\ڰ-�'�v�����?AV@f�\c�\0��C�S(��Pb�|��H[�O�L3��O����O��]�,��l̆{��h`j��s󌄲`�J����(X�����OVLsS�?���ݟ�i5���)<� $��P��	ᵫ�+?{rc�����T�'f��;��cʢa����e�8UB �l�KC�6m�"m�����O�)G�O���'u��O�L���4x��y��*=~� �SpY�iNNQ�'�b�'�bZ��#"����'r^��ig@I�lܝ��DƟ`�j����i�R�]}����?i����>	&��y��'k�92�D�1a������	՟��'*�,[��)���O&���u��Q*Am�)�.d+�&ݗLQ����O� �b�'����O��ϻ?^�h� �7Gs�}��G;� \l�kyrC,"'�6-�E�T�'����<)h�w�-�0���q�x�RTMs&����0@��!2Ц�%���C�|�h��4&ͺ3��$��O�� ď���>��L& �B]�F���<d�&j�K�<���	C� ��4/�=.#����i���ɐ��ѾB�ڌC� �0+�>�!���W�p=��,�32�]rk�΀i�bJ��s���U�1M���NE�|)��˪Q�A���7�<$�H��g��|���?u�L���,��ǖ0�n{g�+Ԥ��Γ�As@�;�lV��?���?��L��q�[���4�I��@�&�5n"���s-L&v"���v�m���#lO� �V=i\̨�B	�x�Q��͋(�m�` �NHĄ�7L5�,��j�����n�>�UBe��O"�d8ړ��'��=��K��u�l��*?^(@ۓX1O"S���S����˛30�� 9��$D���<)��B$��Γ�?q��&$=���6��wЎ�'!��?��OH��"�U��HΧ6���`$[gd �����M�eAP?�n�(o�q�x�� �x8���B���
OUrc֛���mz��G�&E8�'CM"`@| �'O���'��R���Ĭ�rYw�)X�ڬcg'��i��(x K΂�:� #J�/
�	p#&�I��HO�S=x��-�o�3��q���^�VAz3+y�p�'~Ĉ4�<�y��')�U�m�)� X�y��[��@�F���f��Ǎ�O\�$Zl��4�[�m+�	p�O��m �y���3�O�p-R�V(R������w� }3H�x0VBZ�Π�����5���D)
r,ǯ=#��� (f]��>�b����	d�O���эWq��寍�Ѿ9�O9�y��92YV�h����~����K�HO8��S�~�DxR�ܐ�V�	58$e�x#����.SȄJ��'��'�	��P��r�'"P��P�D܌@l9*�J���F@c��\%rP��'x-�奙�k��"?a5���2B�8p/P?6�FU�"^�o(�)J A�7��7�3Qݎ\���L>i&�K+U�>���ے2�� ��-���?�D�i�Ɠ8��,O����2�sp��#ވ��v�̐:'`��!�S�O!�iK/[a��+����&��*�4Nj���9��Hoo��V�SMyr�H�h/�E���=�@��K��ur��d�ҞC��'�R�'�V牬wT�~>�1V��\��H{��@WX�R��X�`N��TmA�%�|�.� u�eo�/��)��C^�ɳR�d���	�X]p�c��+Ԩ�6�E	z/ Rg�O����O\��<�����'�9�MA�G �5#Q����m��E�1O��A�	�1�<�q�M�<�T�s�$��c<���<Q��R%Is���T ��«Ud� kJq���Ο��'I���'X�I� $��0v��Q�xP�bcm�ڌ����; 2^ "vb]/"�����'�F ��B���Jc钖L�i�{�L�"U��,"�P�����+�p<	�ݟ,��ky҄�/o�G�̏F�P�V�B���'P�'n�y���t���p!�b�3�}Ҍ.�S���_��z��������a�ǀ^�8�'�K<�Yz���֟��Iw��@�>�?�Ā�:����3��x
���Ũ�?���4��بSA�����O�t�|�h�&C}�2�� H`F�L;���'w�"<��$R1Y����+�
/�|�D��i�d2h�'	2�'��2a� ��%c�%+v��7ae����d�O���D&ݖ�1%�6_�.mz�P&ۑ�\˛'4i���
Ej,X#G*
�CgZFK�mh���O�����7�z}��-@I�0�T���u`!�D��xI�����=B���+ K̡}'!��]�H�{��$�:9z�O���!�DP��|k�nє� ��׭ņTO!�$�b�P��"�ɖ0��` 7L÷Q�!�D��Z���2��ޙ]�|���IϽ|�!��-�vM�gJ�=�z�S�)���!�D�6u���D�<7��܁��J,�!�� 1i�����]��dE��;$!��
}����"/О�<�q_�%?!�$9�"XR�C�5��Q���  !��)#�ʈrF�A�!����m�-\!�d��c����H:g �9���	�!�ǓZ�4Q��.�+v�h���g�?�!��]�\F�t��,j�*��]?b�!��=m_B!���p�\�95�޽L�!�DA�,�o�Ӫ4��]!3�!��\�?7�����X�P��nʳ�!�$�]�4�s­�� c�q��<z�!�L	3mj�#�Pg��5�����&�!��1{������K�4���++�!�Ȁ;Up�Z4	�1���j�DآaU!�d́l]fa����>�6��S��r�!��@���5`��~@86�3�!�3�Fl���!0n�(�F��2q!��[�"����2���W�ӒbX!�$Q.-ꭡ�*Vc�8���C��N!򤙳zr���f'�=��8xe�gF!�D;wj�a��
�4��ŐbR�K�!�$�"y���D��)���4�!�d�%��1q�[�ze �1���m6!���5L;�r���u�<�a���!�]�PT�i�x�t�
���.i!�D�<p�""�i	�2���0�Z�-d!�D �KQ:`���E�V�d�p�ˀ	�!�� �E��cR�IT��AS�J�<��=�v,_&=66���0��$�퉚P�<X�� qs�;e!�0qZ����=���d�<�Ĵl��=\�iVcQ�[��h����\hC�I9k���:3�#�Pr�ғ��c�p2��ӑ����ƭޯ�H�j��HʊY���ӌ�: �PE`�"O�q2g�/�5�+[-|VX���%{�ٱ2�\A}2����	%z;(�A0D֓k.����@�f"C䉰"�¡ �m�#U^Ɋ'j�:l��(kr*v�n�)]�a{R�:�BTN�u3v����0=i�K��3r����	�~��F.�AH�����(B��a7�Ւ�ykD�lW��;WO��6d��f�J3��'tё�K1�Vd��e=�'{�h����u�A6C��/1E�ȓ)� m��D�68޹˔o�")�� �bӄ�Z�)S�h��!�g~��G����,�!�0�p�D���y�ޠ-���U*U)!P����Cy�-�B�λ]�Bђ4lO��b#�"����Sb��Wʭ��'�V�i��G�/���H�i�ޡ�a�Qr� �Z#��"~>�-�g"O��A�m�-��� ��"a0���W��� e8�Ԣ��Z`�v�F���ƚ)�J��A���@ H8:��ǹ�y�@<c��\a�J!����t�+(F�s&H�r���'�HaE��O���Ԏ[Y��xq1M)H~��: *O��3��G��� �/��u�@��87n�P���ڐ��$D�6�q����<!Fx��6y�Q�L�W)E��~�BI�+�I��O�.��1
z�[p/^#6P]�kD=%�!�DGzpp)�ݿ~jf��1�tT� �VqO?���g�^��OW8-�� �2HV��!��4o鈐#޿%��`yAL�G������D>Ei��ݦ%�2�N. ��ɪ>�h@ �O���&�-�!;�ΐZ�:��'�j�䈌�>�#'1NX,P�B	��d�*���t�-`�OB�P�����K�UKfC�	^ʉ+��_O�lU+F�̅^V��`���f�OF�}�Jff�H3�xL���Pg��h�ȓ$_�s�
"&3F�P����"b>��	2�  "�c�O�`�C�ќ`ar�r��.F�`ro>|OhШ�d"���I.D�K��.R�^`I�=%��C�ɾ��q��/X|R��u��$�b��V�yP)D��/� r�5���Ye��0AM� �y�a��Q:@ s���|�n�Ǖ�q�X%0���h���n���:Pա;O�-�Rc��+�!�$ֺCT0=�%F1OB%šև1V�ұYr4���'dB���8�X٪�۱~#
m:�'��@"Ʉ3�Fd�f֯q�q
�'3N�4k�	c������>i���
�'h8����ZX�Y����f�����P� ���S�{���fZQK��B���B�ę��=	 �"0B���D�':�0[�L��L�2��@脁.�<$X�'����M��1���&:d�����6=�!�,ڧr@��XU	��R�@���j=�5�ȓC�9��D�C�t����&n�
�x*���Z$y4�>���O�����U�Z���V�]I��E��"O���p#F�4�2�&��6&m�����'?r#)��m��L���8%���s �vn�!£�U�]���D 8�J囵i�:�Msf�V�h�th�/7a4M�S.��<�Sj^fh�I2�E����&��}����������̚6�r	N�'����A��4Ys�}��9j���I�$<�DYקƻv�PH�.��>MU	'#8O�@%AV�l��53P]�T��JG/B�H=x[H��#��o�(�O\�ʓ�'r���5 �&�tL���40�TI)O0�5E�P�!*V-��~<>��S���� ���TC����m�$� )�ȓ ڕ�qg�	I��lhG��h���	�M)Z�6��شMmH���G��j��Ϥ��OJ<��K�&��iytcW�9��w�!�O�5zRP7RE����QP�T�1/&}WV�"Q�I�Z�C��[]sqOҁ�f�"�)� v̐��ҭz�Dmpfo���k���7���ɉ�!^= D�A�]��8��d�<��!���S�x��� i�i��Z`�'=��Ѡ�I���ց�D}���O`t��-Y�J���0s���!&��4��7N�B�.x�F�yFK�8 w.�zt"ORЃ"�!�"���LU�.��ũE, }����#>MT��M�D�)�#���d_2�n�C���B��a
/�rB�ɞl�ڐ�qd�!x���E�ߍ~�4՚�+X����HD���c@CMx��I1+�6W6���ŀ�� �� K:O����m�k���B�%Rޥ�·�5��y����z9bt��7y�|C�ɰ~2���]r����\�@z`�vd��S��2���GS&;��m:�S�/Z�DhF�_h��<�v��zd`C��1}�}�� *�L�DI�=ք�s��7;M "�J{Ӕ	+2ϋŖI��'�(����W(8OE�B�B�Z�>Q��'(����@B�̠�R�`B|E���1�5bp��,Z�(�
"�Gh��R|i���d��r�jt9e�Y�ў���O:E�"0 ��Z�NXpR���p���G�u�܀ ���I*W�'��x��2,�,R�ԧSjZL˶�Ƀ�?����a�L|8��Ք,��=Z��R?��i�f�@1"`�X�kI��yFÈAA�p*�.S�<mZ%�R-L�}�4�L��?���'U�u�˟�dh�{B�A4 �\P���
q�*�&���0?QL�!�?'*;8�( �uB�(D�aScߵ1"���ǆ2��pD,,\Oh�KV�!	��@b��\��)����d��]0L�6���B�h�IRf[�.��}9���-���� !��$��;ClԂN�N���X1_�1ON���H#�B����(�ʥS��A�~[旂\՚�ضK%�y2L� @�h�!3��g^]JFA֟_CD	 ��V?r����J2��D��OĹKb�Q?_�0q���a��`�
O�$�k��TqB�̑=�l���	�0� �@$L����Ol����4t�%�E�_|bT1��M�(ax���������<�"E+TÕ"40:<�nЌ&�2)Yc��>XxQr��c(<ia0V�dزW@ՙT�0����I~b���s)�`
7��?R"� ��,�?9��4{�0���A@/4�P���	�8 HB�	7 ᴀ��hR����ʛ�_�qF�k��#�a�O�ظ��u�S	@)���!�a�E;��$��H�5��?0�����?�D9�R:�舘�$�:������^�+��#P��ʟ��7�
�}��d��@^FM艚�,3��+G����By�g��,$��I<4��[��)�b)A�,�֝/A�d@J�
/GԴ��ue���u�C�]����U��p:�o�7�4���kѐ�+�f1}Rc�_V� �SF�'����.��?��%��y��
��%�t�,)�v�K��߮{v��ȓBP�	27�R�w�LD�� ��+\hZ��f!Л<����<�O����$�k�ǈT�!�/ұJ���KAH<1&�>C���(���9*��	b�'��qP��S����o�5`��}��E���}B5�@.���5&�/��<A1�P<n��1.�^�DdՎ1�ƭ �U4R�̕��)�9E�V�f�* �\D!��Ly��P:�GŰ%�<(�)��.�<�	��0�ɪnY<��� �s�TY��ݣ�OT��#ةB�vH�4���	(ɻ�b0D��Se,I�e�� �ݛ� r�$TF�Z���.�м���@�)��	��y"^�wnX5*�N	�q���P��X��y�j�e9p����N
%sJPk�n��V��'�敢��̀��Ւ\�t���*��S�D���"Hv^�R7�X�$�����E5S��H& �:O���pҎ�
y�摘P)H�L���/gm����g�Ia���'{>=��l ���P�D	]�E�6}���`ǆ/��}x��� ZF����������?L�E������"Ov��2�\9�RH�F�*&|A��o�lCΔ�T �$+��`�O�i}��9��1����6����N��@$�"O�)���ř@�n�����O"�&F��k^\�I�;z���,� (���\ *7�O^���`ƾO"�S4�Ѹ1ǒ��3�'�$�so�+WRA�֣��H�>ـboCP�%����.�J����-hv6U��ɋ*� �'�	�^�!Ku��.	L�=1��چA���sF�ǙHR��CS"���$��졢��2BF�y�v) �y"�|����d��J�V@��!��y"aY:�(Ѩ�ed��!xz r%
#`��!	U",H�C�?ђ0Y�G�� �|�j��'�O��x�������D҃��)����B�X�x�!��5M�� L�"ef� F��35 *0���MH<�d[6x��@F�a�TXQH�h�<�%�$w���&��.4
�ky�<Q�K�:%ܸ�P&�]E^��
]�<y�� �N-��D�I,��wH]�<��c�^n(���j�=j�d�DDq�<��JW�e:�*F�b��dh��Yb�<�p����M�e �;�H�֡�R�<AB��mbл��F�L(%&FR�<AcƩT|���]^�֙[�(�Q�<�U�Į
�蜐3�f�HcuL^J�<I����d��=�?V[�3D�F�<��9I��4��;X?R1`q�I^�<!5N�?2�Ds�'ѵ\l�F^�<�G��$+�P��@�1S�ze۰�Ls�<�����3�	߃����eXI�<�C��(S����XK DC�a�M�<y2䖂\:���ՠR�y��R�m�Q�<�T�`+<�@���4G%*hQJ�<�.O����a�������W��E�<��r�ٳ�Z�Ն]	!�B�<�u��>=��r�!S�d+<��5MJ|�<qS�e���Bq���UD��ā|�<�G)F	 p\��F,s6ؑ�J�y�<y��$F��-�Pkǩ�> �̂p�<�����k.�u�'��H�0Xj[X�<��
l�j��6)��6�xp�G�M�<A�%̝x�Re+R$�J����-F�<�1 1=��:҉F�*6�U�"L�<��e
�T�lUy7n �b�Q��^�<!c+�?&"���؊Cڂ�S�N �<�r��� Q��-�5�M��S{�<iwL�'rza�Wh\;4�Ͱ��l�<i'Ŏ�*ǘ=*w��S5(�X�it�<�� Ϻ��Xc$�E
<G~1b�&^t�<��iJt.d@��Y�
���$Mm�<i��[�[P,퐴͎���7�]t�<�^2H��)Z�N؃P�����k�<	4n�A�)26�>U3�AT�Zk�<��Q�5L��V�9�~�� �j�<91 [�y�P�U�ߏ	z�%��A�<9T��&Z�Rlp��A��r�NNE�<aa���/�ݠD��6��r��|�<��#��w����ɕ3��4�a�<ɐE�jZ�4ҌɎ)���"	�C�<Ir��R�4`��Dİf��q���P}�<��#E�KFN�X�I�+��!D�Lz�<�R�"gH��$�ة"5��G��w�<Q�
�;�0xA��V�R9�Vp�<�,��}�,�x%Or��`W�Me�<���7�h��MA��ms��`�<�Ύ-O y��F�k�����]�<Y�G�X�\������+3h��t�Y�<96�ǎu��`d��;�v�A��V�<A���_��,���.2�\�vo�T�<Y�fd8�03�Ϫa��McG��L�<�ר97��]A Ü�Q�5��n�<q2��	h �H�r��%��C�<A�$O�U�&lj�Mɿ
�0�bQ��{�<13M�b̸�����&������n�<���ʇs{�9p)ѽ^�U��Ãh�<i�.��"�����Y�v���L�f�<��A�~�����n��)�R�!�`�I�<�f��?)��ٗ�T�<x�<a��D�<� `����7x�R`ie�'B��P"OIYsj�?�V�Ǯ�qJV8x!"O���C��94�`�+e�ŉ'N�m��"OP@���4��85��W36]� "O�T9�.2��)pbjO�q����"OvPg�F#yS"�X��H�6��k`"O�EcA�<NT��nG\4���C"O�qm]`p�_1-���"O�I�hAg�d���3f�>0�u"OL�y�I'l݀T0^�0`[Q"O|ى3,þ;c�m�SJ�Ţ�� "Or݃�͕FD�8d��OJ�B�"O
l��$��.��(6c�T4��"O���ʍ�?SD�@%ŷ;|"XB "O�UI�%%*HX�2$�)y�L�"O����*�
r�%����la�x �"O���/� ����@�'VZvԡ�"O@�:WkH!*��<��`��عu"O�2��>xh1rVFǷ��DC��,G{��iO#�<M�ӡմs1$|1§Y�9���dȿ8��\�g �sb�cC��7�yb�UShd"�OA	��Գ��y®Y��Dq���d)���ֶ�yR끄(&rxC��fI
ȀJߍ�y�c��x{��a�p�єB�;�y�H�*b~�Mh☽���Ȥ��y�w��z$^� <��h��%��	|���Og80�ԫ%3��Y"��)kʡ)�'gD��WdY�S+vDY��fM(K�',Z�b7�һ5���am0ch&�C�'�6h�D(-Wq��s��H<bV\�'�%�+ñH$�D����i��'ɸ�۱�&@�Ba�'oÐz����'�-+c,�#!4���)-k��9�'�R���X6%�Y�f 	�8���'lUH��C"j��4(�߹7U��0�'�X|1F��-b`"g0bҤ
�'��	��ݰu(�0�@a]I��'�&-�%��"p4�
7���SF`��'��i��b0�c�`�7� �{�'Ӳ-��X-����c�JM��';���M�T�v]X� ݟP���Y�'����JդqS�QcJT0�P�'�d8@r-�,6�"����Y�P�	�'y�xig�ض5J�[s��K��H:
�'VI7�ݔ"1�Y#��7O},�	�'PU�s	�������#@J���
�'���t��/dB`X��D�8��Ui�'���KMV�
�x0� �Ve.qI�'�HKQ$@+q��T�&�M�DM�'��!.PJe.0�u��4~P(�A�'X�`�CM!D�%ڢ��"@�U�
�'B����/o�(�hU�I''�h<B
�'�}��&�}�|��t��8��L3
�'�(�3�سW������Ė���	�'����$�+�0�E�P��'�E�g�	�B���	�����贉�'+��9T�Ґj�Ȝ�B ٵ~&����'�ꠓ#[�ii(9P����p^�iP�'A��3�h[4i��c��1 �|=��'�vp�B��#dZ��$%Y����,<D���soC�k�t���Ҏ%a&�%ɾ��F{��I�r1� ��N$�a� '[�!�$7n�r�8�B��k�|� �֯; !�� ���ʖ�a�x�c"�v�`	�"O�LY���!@�h0�K�rK���C"O�����B��5 PK]++���"O�E��\n�P%���w@Y�$"Oz�ǀP�P��Ł�D��, "O��x�&:w��5M��|d�!��$|O�$��lПAl`Yfǀ|��3�"O�ZT)U:I����D�Quq�i"O�\Z���T�d��`@#_]ba1q"Ot$� 9�A%y)�{!"OB]�"�T�����J6�t7b$D����/�* ��yvOL�sh��5$D�0Bf���=�Z�(�]��C�� D��+D�(R�=�%+�fH�����?D� ���R�J�v�I��ZLĀ�7b<D��`s�]�9��-a�)&X8�`S�;D���䂗��I��D�R���Zֈ-D��Q�M�7�D�#�F$1��XA��>D�H�5)�J��s �<}��Xᅠ<D�̨�kƀ7�<�	�bŵ|=��R��;D���ּM yBS��<K!�I�%o5D�@k�$L�r����l�,/R9�C0D�8K�F�t$션�'�m(F��0D�x��� �bAi�N�0}.}�'�"D��pA[9���H�N�N��)?D�d�@	\S�P��ӠH�2.F���)D�h�䀏�/w<�r�)��=k�'D�`�2a�'M�9�k͐o���P$D� Y0*��Hj�B���,<ȉ�׀#D���%���JH�i�ス����'�4D���RʁHD<��'��Q9�m��i3D��[�(@�NE
�_m��h��1D�싡!u.*Ւ�" C�m�@c/D��) ��-�|D�À�V����2D���5*C�̔yp��!���P��/D�$�	9t!J�ŀ�{ܥr#
/D����C� R�ڴx�Mʢ2_�E���-D��1��S,hq�t��C�Q�Rڇ�*D��2�T�gB��!���#� �z��'D������4��i{ �M�K��0(��%�O��I�}�����F�a^�@���U`C�I����P�Q�,����W��X�>���&�Z91�̗�u�}A��:<�>C��m�N����K�p��`���$C�	�U�9����4"�����A��B�ɔ"�б"H�)LN�2�H.\NB�� i��H�UɆ�@��\C��2;B��3��%p�ϗa�P�WQ�V�C�	7c�v�����@Hn�i��TecC�	l^*z!�ȪM�F8SscM(50�B�<�����қL%�pGō�JzC�3Udy��>U�$҆�	zbC�I�#�d-���a�`�[Q��!QRC�	G���k��.l��ȃ-UBC�I����y0��!6\T��S�+PC�"?Nfee�ם^��Ԙt�֤[�B�I�,��#º0���4�:8�B��4���� �e_�T:	E)��C�U�>8��b�6'ټE	�̏���C�	$q.����ם��(�'9�<B�I��"F�S45-���aO�7 B�ɻNM�vl��#�����,�C�ɠ.�l��JI��n�"���B䉬cv�2�nݪq�p�%�ڊ���� ���,D�J��-�j��(���	`"O�ïɚw"�.չm����P"O
�[W-�10�zU��$@��A��"OT��T�nW�ek�&��[I�h"O� ��>v�� �#��H��ʥ"OЉ���QbJt 󏈋fѺr"O`���Rx�2�aA \f�	2"Ol��nA�L� ��vA�4	���"OJ�6�FU�@�%��v��"O�i�&ۑG�<8� TDcfq#�"O0�r}�BPf��`*�=��"Ohy�!C2:�օ0uC@�K��찠"Ob|bF	.�n�0��[�W�Z�!"O��K�$܌-��B�8�*��b"O�i�����J��%�!V�8�֕"O�p%�מ%��a�/
E�.9aV"O�X�3�2"R!ɯV��e�A"On=��Sx�(Q�\x|��"O�Q*W�"X}���T-�;<q�Q�W"O�	A���RiABL\�&Rr�A�"O �j����sy��(E	��gOL�q'"O4ma�g[�As�0� n>nP�B�"O"	CR�I)U��}��m�-\�c"O�h��H���|r�`^��7"O�jC��!��6 ��KhfE��"OP��QK�0Q�]3�
� ]���"OP��AE�|ʴt�W)W(LP�,QU"O�E8��=b��a�nI�;ޕQ5"O��rb�M�:��0 "n^�IS��2"O�P��F�~R�!2�MީR\��"O�����hr�L��B<i�e"O~V!h��'(R�z�H��� �C�<�E�S595�M�MԲl��E�<�e[3-�T�'+Ld�`��h�x�<�����230���X�"g�=0t��y�<�thO A-��:0mZ2	xQ@�y�<Y��O�Ah��5�B�L��Sw*�\�<Qw�V F�4sp�Ђ(�}�4MH]�<���ˊp� 9��ӺS�0��憇[�<��!D?�^��(�8#�6�z�l�<T��p���x�̚ 5@yZ4�e�<14D��TH�#[K��!gbZL�<��uI)x��ߧY
�VF�<� a�$������G���$x�E�E�<х@�)g�J�!me�1y�k�D�<yT�B�D�,0�@T�*]˦�F}�<�q'�!	�EA`ξn@��*)Q�<��&��u9̜�J�2l�a��P�<�0��ck�aI�B�'Y� ����U�<Ic��'�
���!9�0���J�R�<po���>�����
�xH9%�J�<��薪:,>���+�3����F�<�g@��n#J}��	�e�윐5 �k�<!e��%=���F'��0�DP�&�j�<���R�|�XZu�]!�L88S��M�<q��\��ٓG� ����HEU�<�O0� Kf���-Ae�CN�<�GT�d�2H���N""o�e��eUI�<��)��6O�e(�(�����##@~�<��}8�`$�
���@�y�<1R��/��(�a4/�V  �!w�<����9����瘳x��4bd�r�<�W��]�����HƵi�>��Fl�<����F�j ���߮��9����d�<� r��O�25�$l"��=Mu.!1�"O�i���0��E�t[P��"Ohp�,\�����J�&V��Z�"Ov��o ����/�Z�j"O��)�͙(�p�I�E֪��c"O����I�/a�\m����)�p�i6"O�a��Ð<\��f$�"Fs,[�"O�x�&��Q}t�YQ�
a^��A�"O:!�i�21kL���c	J��e"O�4��(�	?T�P��GR��"Odٰ��U�w���'�Xa��Jv"O�TA��7a�t�c H�v
乱"O�;w%�"}��c�/ȱE����"O�Q�2cH'��H:O�-1E�I�u"O��+4���������dZ���"O�Ͳk�+X��� ��&EV���E"Oz���h�:qs���l��2A^���"OZ\�tN�Q(��y0K��^;�x��"O�����m,�X���2�J�"O`�P�Hǥkм-���S:���YP"OJ݂t�1O�$Q�S�ݖ�6Y�"O)qЯ,��%���5"O�8�h�?K�z��#1j�eHr"O�!)����r����3EʥVg����"O�C�h�82���u#�4=g��)�"O�Ș$"�%������V1H��1�"O��xbAԢ�$��� CZ�+"O(�A&�[��C��O���"O6�:so�(N2	2�n��p���$"O�Da�˓�u`z���p���"O�8�KCn����Ջ�'e�����"O�5�e�T�l�X�`��P��x�y"O��l��*B �*�iP&��,�7"O��'�W�(5�P��i�4'��d�@"O ��d�9�V,�B)J�
��Hh�"O2I�$�i����G��t�2"O��7"F�u�����gC�(h`�"OnH���D�:ܛ�F���|0�"OPh��/O'cq�*�%�+���'"O����g�+gf�إ���az��b�"O(��7-���������s^�s"O��2�R!((���֕Y?~8{�"O�
�M�;|��C/�p1n �C"O��a!d�,f��i��
>_�a '"O�X$ψ�7,�jց�F"O����jI�K��`�G����4|h�"O~��'�âj�nzd	��1+�<��"O�|CФ�#x�<X�oI�Cf��5"O2���oR�!)��� �1u<[�"O6j�A؋5��0W�
<E��	(�"O� ��V��=��ǧg��`"O��!�o�~�Y��T<5��"O��I�A��&gH�Z�Z����� "O�-"�k��m�(�P�-іL;�"O��Z�-Ն7�}���ОJ��y�"O^@��)��*���aX�Q��A�&"O�i��-�2�dh�؞+�����"O�M�a��yrh�r��-p� +�"Op1#AY9Hf���Ȝ�K4���!"OԑA��� f]v�3�(P�Ԋ�Q�"OL�IR/Ĩ,ifa��D߄-ˮ��"O��	�&X�s� N�-+�"O��+�	'R��p��eB���"Ol��hX�Ԗ,�w��&H�P("O� ���`l�-��#%3L!�ћ1"Oˆ�F��,�1�4�P��"O������c�,�W��&�\���"O�W�r��1m�5����gm�a�<)�	2�4�:�ʆK���F!a�<��j�P�f��4E�^���tŗ_�<��	0�ԙ�����YP����G_�<!ȁ�����ը�z	�.�\�<9�Ԗo�,��_��
%�#�r�<��jK�)��4R�ʅ�5Dv���q�<C'(5i��I+�&DAOVp�<	"н!��)ˡ�N����k�<ɰm�8S*	�I��0�i�ŉg�<)Eʆr/n)��ˎ-�U�be�<	v�����UEh\�\�Nbƍ��-0�3WGT�(m��@�$/����0��$(ELœ|%8�v��ɔ܆ȓ;�\ˀ��#�a��� �.��NaT�����nȀ5�a�Ƒ ��m�ȓVK���+�3?�����iw��K
�'t����h̍c5@���I�&{�r���'�L�Xs�9��-	���:m!Ȝs	�'h�葷�T'R��<s�J�w��e��'d�"��%��y��]�����'S�q�ₒ��`r�-MWkx\��'a���#��-z�l�0�$NF8x��'j�J�jا�Ȩ;�@&B*�)��'���R��>H�(}P��QQ�@Z�'��-��(�! MФ��L�:i��y�'�x�ۂO
�_CJ0j�
,��8s�'t�����Xg���Ŕ/9��'o~=�d̆@c��rv�����G�1D�(2րT>,b����
!̴ٗ�5D�h�DO&��9��V9c�����4D�Ѐ��b�^�AF�>>t��H2D�HPD#i��%M�2y��3�*O&����B��`�YZ>h�"O^(sТ�\�`Q��x2 3�"O����y��'�Ӵc��Ӑ"O��6L78CvH�� x�t"O2m�b��d�60+�l֥?p�|""O522F��C<́��GR���'"O����4=O\��,��m=�9�'I�I�����&�Zy��#�{ �''a~�%��0��U��
K�8p�WL�yR�W^#*d ��0!�P����;�yRFH�Aj���N�%Q�)�f��y��%,��ͻ�D?N*���ME��y�(-,`��7��8����`���y"/�|PD$"W�_<0Dy�7���xR��b/�  �V&��p'IJL2��ݟ��<e��)d��`ċQ�2z��7��N�<����43J����̴������TG�<Y#J:�zCUiM+[�~�b�+]A�<�eD)�@ �<\�V��nO{�<��D�9�:}
�i԰y�Pe�'T}�< �Z�[�����[�X�l!"���v�<9p,�S�E��N��
����ITʟ���r��?���?��O �a�hB�P^�����9y�.�JV"O�l:al�(f��ȉ�U���!!��)�fqsf#K8.q�i�/D�J�!�DƏ\4�p�H�r� �V�)\�!��٪<e]YF[�8�LB ��M!�_.���h�+��A����❚��d9� ")�fiߖ�:@(ͺM��kR�'��O���0��e�q��t j�I$'�>D���ȓc�0���ԏt<i��O�=�FЅ�u�~l8U�]�W� ��F���?�H�ȓ1���	`����@��N�LR�\��=�h�$�����C���-��q�ȓ(׎4iG]:c����6k	����ȓW�B�sÁ��]!h���0�n!�Ib�����]!4eF�Y���CfB�H�Ќ���5D������6��Qa4��M���B�I�O��=E����`\�U��/R_)����k�~b�OR�=��ҁC��M	�:ѧ@WH&D0�"O�|�P�\�Hz���w��`7�|;�"O�)�V'ܮ&�@��`��
	zȘ3"O�Λ,����C/��7몸��"O E�s��4d�l�;��@��:Di�"O��h���&z�Fa`�R5ր�`�"O�Ti1�ɞx8V�E�X0 �0�|"T�\�� j#PA�CK�>]�t���%Ăr^B�	20H�AץQ�>�pX��=XB�IP�����HN$bL`��ζ{B��4	��	8W��k�~����߁U��C�	�=�qSPK�'N_v�� ��!78�C��9H:���O��:�fd"�k�v�\C�	�A�yȰ�� �&�В��4$<8㟠D{J?���m��p�"���_/~��	�1D�����ee	2.J�#ؑ�C.D��v�I	iNBq��'L0�EC�,D��y�&�0Ub��寚
5�a��@+D��ɖ/�,<�t�T2F��ћ�B)D��85d�g�P@�f�+Mt>�
6�&4��
E�Md��pc��2/N�u
T�'Fa�TO%,��Y!�v�45��,S��y")�Q��IѤ#_ha�7���y�#ԧ`Rr9�b�\���B W��y��6nŮ�QBʚEˠ))��2�y"�L�XP��9-�jЁ�����$�OX��F�Sg�R�V��
C��թs�'�bg�P!�q��d��V���(Z�!��y��rӢ�=7Rj���ͣpg!�$�$����Y�Q��cA�N?oL!�Dp����r���0Nh%��H��8H!�;4뼭	��M�G!|�c�g$�)�uE�<{c-"D~�� k  /Z\p �'w�#0�I)lVT� ��vL���'���ʅ�~&$�H���?/t��L>����0=���֫Y⮄�q�F:Ab�s�@Ra�<���C�ꑪ��ԾB�&�J���T�<'�ڎ`�ѣx>ڀ�$^�iR!�DYr��ui��Q}. ���}T�'Kў�>=����dU谁L�D�z��A�)D��{v��� ��g�&>a��fh'D�|�')	3�����Fd�ע�<9+O��=��B��r��,�2�;>����"O����ɿ=l�����6A>rѣ�"O>�`ԈM�m*0₨�lRm`pQ�$�'@ɧ(���9�ŎaCJ��ugٯv��"Oݻ�̅zR�x�&[�[����"O�Y�C�H8��dՐZ�D�0"O0SP#��Qo`[�C���`�|��'�xl�2CԌ	��!�^	f�&
�'\İ l�.�>C�&��,��'�����D�V!�=�����-�u�����$&�����u9%�°l!�I!�PK`�	��S�? �}��K�.u
.�d�ۊ��"OB�#�݁XQ &B�3�t"O0)ВΚ�8���A�eTX�x��d,LO"ī3l���b`D�<����"O2�)��G�Xz���"�٫ϒ��u"O��en��Y�!-�&��0�"O�E��� ~B!���B�L1�"OU�2�Oy���rc�����[�"Ox '�(!/���q"0yx��ط"OT���Q<`AX��R�,Ԫ�"O�<��(�J9�5�#�ٮdKnE�"OV5��-���� P�B������"OȰ�R��^M�����đv�B\��"O��pm�|H��$^%V�p�"O
Akg�1n1V�q�cM�pY`�"O����B %~vɺF"�7u����'$ў"~�-�1^�|c�j��`p�4%���yrO��i"@	qp�U'84B]ѳe��y�R4�\�Cc�]�$88i3N/�y�C>�x�%ǀ'���;f�ӽ�y�M�4\�hPB
A�Lf@ɒ��G��yi�~!DZI��I��)�y�/R�zO���% �)t}��`�oQ�hO6����0�8=[%k^�q��чؙ:�!�$�%>��A�4��$a}:�*��2�!򤌸�\T
c�m���l��=�!�bb`���]#u`��Ǭ�-1�!�Y�2RH���O3R��s�`^�џH��k�Oό��C�^�H�Jy3�IA,Fd�bߓ�?a�O4A@Hˎ��X�u���<��D�s�$;LO���D�O	�8 ���`�x��	{>Be&3����@��lF��u�"D�l��)Y3f|pZ��ύcLLǅ>D���O��M4v��[��pӈ\��y��WE�@�Ӄ^02��������y�_�%lH2���?>�P��ĕ��<!��?��O� ���̒��}����<GD2����|��'qL��@m�U�P������`�A�'&v	�a}~j)�bb�2e��#
�'��ҷ˟</�:iY�g��1�J�	�'�J�zG�>u���k�P��	�'�zk��N�nt��C�>(���'v�� uc�;m֘�x!Nľf��]K	��?	���y�@��b1$�ZQF���!ϓ'�y2H�0~�X0`!�:>~�d�ԉ�yr���s��U��/<ݔ�z#Ȃ��yg�'������]�)��D�B���yRo�F2����)���+Q�D6�yRLC.X�Y�(�(��X0����1�ĩ<y���v�P���+V`�0h�a�@c"�)�D~��	o�4�"�ܞ!N�]�0�[��y��
�;�,���zL���!��yª�3F�le�gؚ?����yBfC����pecd��YEC��y�HP4.��-�g�ʯ	N4��+���yR�Yb��Ȼf���n� | n֛�?1���?y�<w��/�8MZ�5/trm�Q�T]�<1�kA_��c�E�C���fL^Y�<��j��4Nv�x��G�W�f��c	�U�<ᖀ� t.tI�+s�:`�"fX�<1g�J
E�M�ӭ�##:�	�S�<���=�t-��I�Q��(��`�T�<	TK
�lL-�p ɖ+�@����q���?9�ҝ� �à�~�x��cE�**�(��9D�� ��`�=y^m���>n0s�"O.�ن.1�
�+g	B68Đ"O�%�Y�y��!�n�&F�h��"O�9��#O0bƄr��Ҝ2��k�"O��W�KPR�v�Z4;zTp%"O*%Z�W?Il~l�A�&oZ8�X�P�T�'����~zWA�����CY>"�H��ċI�<A�m_�.g��Ǧ{s���P�E�<y��F,; Q�D��6Oe(VGBv�<)�W�^�TyPĢ��-/�h�@��i�<)׭�:\�4�D�4��ݫ��a�<1��J�o�.A �&P"��S���s�<�&�!p;]�c��*GU�t˓�Sn�<Q��
;5f����R HJ��p��q�<����)|0���gB<]�FU�$��h�<�6fE1\�� @'�L��h�a�`�<YqM�,�nl[�+X�����W�<���	!\KdxcE͏r�h)M�h�<�q�ؐ�~�#�_�t����W�GO�<�!EP� �4���CU�UUQ��/ß�$���	L�g�D˹UnE��D?
�t$�B@�%�!��	o/�cB��w��M �^�%N!򄍳q*��9#c�8W�,�Ph��j2�)�'�ލ9����Aj:0��E�8��(��'FV9'j��<-����+�`�=��'�y�"�U/���$�P��ܘ�'�@�Kq眵4�zD�#�!�"��������>!� �zT���aC�|������W�<����$``"��"�S�p-��;�N	n�<��%�=�LDXE� �s��c�f矘��^�S�O
\{�'�>���f����L��"OP(�ĬB�+�p�镡1f��4B�"O��a" �):�u�&j��D}\�x"O����&DQ��)������Z�	k̓SM6Q1��;���cƊX���ȓl�}h"��-2�QSa���,9D�ܐS���&7��k�/4GUl��Ue�<��哆G:������6U�(��� 0K�B�I�R� !�1�ާ:=\Y����o'D�\�^�+NE�b�;Լ�*�E&D�xk�:0���oR��� �!ړ��ј'���CQ�%��s!n#zXH8A
�''�Ҭ�)u��E��+7ti�a ���'�a�D�E�i!��*Ǫ�WɄ�9'%P��yRą�#f�Uc�^1L��@	w�F��yr�Q�+Y< �`R&@�(�c��̇�y�/��1�pĪ�Fťs
|�u,;�y���t�t\H� ��h'Hf��)��O��$'§P~�0wfN�7E,%{�C�0�\���~�z������eX��:Ƨž<H�?�+O�#~��i e�E0�+��4+� �b�<q �QP�c�˹2\�A%�_�<�];���S�&�0Y&���H�E�<����L��f�x�����C�<�*�P���'�:�r�1��y�<��M��iIĬJ�i�z���K�<����Q�Xr���� ;��WG���?������D�*W"�sv.���DŮ'�>���'�a�b�ޕP+�I��/΁�2 H�'���:#:J m��F`����'�� �7~v
q`e��map	�'f6p�����	2C��]n6<B�'��yi��2^�T��5"s�%��'��aB��U�F$��� �b�jM���� �9@��56�H��ԯV���F"OƩ!��G�P�Ȉ�U̟�i��9�"O.���K k� 8��*&o��B"O�ŌԬh�z��-7a�Mh�"O��ҁBSpU�"bΒ�q�z|��"O2�b-�1D��H�ƫS���dYs"O��{Q�aކ���g]W�z8iP"O�� e��g�u�4���#��K "OF����uR��eQ�L6�@�'"On�6L�
0U���Şl����"OTM
Ge!;ĺ��_�hd����"OVLR���G�pBN �EJ�-s�"O����I� �v�{�@�[�7"O8sb��*M��#��g,`�"O}#��beD"�!AeN���"O\UBq)�`>:4��͎(}*Baʆ"O�q�� ~\��p���t�!�]�el�����UL`PQ��f<v	!�d��>/l���}R�3�c͡O�!���V>�uCa��Q��|�R�۬�!��%�DZ�f���KF�8f!�d9?�U�����n⎵�ѣ
�1d!��'[�!�d!��N��؛3C1]�!�O�{ ^5X#�Z9h��@s�
�T�!�Đ A'JᐡLG��I����!��,w���Z�J�?a4���o�!�K�s�䱩p$�i>1� ��]!��E�<��T���I
rxb9���ԯ3ޡ�d�V��U!��&��a���%��C�3d ����~��rF�~��B�=D_��Ji����!�h����B�I�=@\S��#��,H�� `3C䉣{���H���ln҅Y�H�sy�B�	�=l�)�Dd��x�v��8;�B�	��J����y����G�MYBpC�ɘK��u�$*D;,��8b'λ3�@C�I�*p	����m"�4��(��i�@C䉶u�nžy�V�Qm�?W&C�ɏoG��Eʗ�QT�Bgn�%`HC��.rmYg,	V&0����\$��C�	;%dD���NK�J��&(�m�C�I�\��qwb��W�%�`�R+EڤC㉿\�h�� ��lV2d dA
t�ȓ/��ԁ��
�	���x����.CҨ��)	�7���Α�<� P�ȓ�@rtg�w�R�PB��U��#;x���a�U���0�'x�d���s���G�T	Zo�h���!3:a�ȓ9�$(IB��F1��ktGY�O�6h��|�\`qR67�V,�%/�*w�!��a<i�͚Gqx�� �Ӷ�D]���L�<9Ѕ��N��`P(�4f`����p�<���X�i�"�ENhdz�+�m�����O""|���ߟc|v��(�T�Sv�D�<y�Jə?��YCK�M`DC!��Z�<�5`�+>nN0ё��a���p�'�Y�<!��[)�2�Y�G� �BiȰKS�<)5$
0s�����K�@�x�UP�<q3NL�=U\ZB�- �^��ůRU�<�6)N*4K�H�0�^�XD��M��?Q���?�����EA.@P�mI'K��`�&�H�C'!�$P�8�A��BH-���K�ri!��8�e� ��:+1�!HB'� Oi!��͈;���-Īa��P��`!��  ()�+�.xHvL���.6^�I�"O��ܶ5d��gh�
`��"O��#P��t�@H�'F�-Zw��_y��8<U]�GJ)���!��??C䉠E�@�	���FiX7�
��B�-u��� �kP�i�Z��ć�1�C�	=`�,�p$������B��C䉟i��,��(�$i��E�d��B�	�9J���p�R]�6�B2?��B�	�xR0h�g�i�Ī�A���G{J?� 4'�
	0����ތg(���3D��ǃ��Y������@�.tP�<D����N.J0���ϙg�,��!<�������EF��QZ(D�Z�(U�"O��ڢ�ڡ�Y��g	*�<:�"O���2�@�:H �[�l�v��"O���i��)��4/Q�U �2"O�Mq���3Jn ��3o@YcE�'~ў"~Z iP�!�:p��NO�s{�y�ԓ�y�����(>f?R����^=�hO����O�"|��;^hn���ˋ"Z����i�<Ag��C��	j�RJw�q�d�<A���7s]���-�n}�u�~!���vm~����qG^�@aA\Pn!�d�(^�Z���I�&g

�S�.Z)2�*�g?AW ��l���bT�S'v}(<�@iO�<A!I�R�}�G��l+6I���r�<�A��+�aC���`X�$m�<q���%��i�鎟x�re�d�<����7�f��'��*��A���K�<q�O։[r>h��� 8MPE��l�<1�A�>�Fڢg�%
�bNB��4�?����O����
��J��ճ��@�q8Q"O�Drb�/p��	wJ�%0���"O^�B��:L�� G�+s#0��"O^ɢ���Ok��#F�
+!��`�"O�9����"=������` �y93"OZ̢"�v�=�"� e��X�"O���Te[
��!I���&"O���ƪ��N�X�Ah�{�f�Aq"O`R	�Q�&�Q�(X%���Bv"OXL�0��'�Tp��#�r��"OB�;feZ�%�e��J�u�"O��1h�$��t�I�	(���s�"O�`A���A|`5��'د�P1�"OԈ�+ƦAh�����9K�>���"O�82��FR�T)\�r��A�'\!�d\a�|���ͧU}�7nG@�!��,�VP����+�8�tB�|e!�Dȡ#�� ����R]�՚�˖�KW!�DG3+�j��7@�Th%�JԇBo!��'w���G� 5#:��e�X�S!�D�5h(<D:4���r�p��V�V?!���:�BYhvA§t�`�:�MR	77!�$���.��7`ޒ,W�E��NO	`!!�P% �PE1(��\H蘃P-�>�!�$�(&�<R�����x�c,�/�!�Ā	K�=6�ټ>[@yx4nکl�!����m��A �	@�M� m�- �!�D���2��a�أ1���!�;�!�dֺE�H$�a��=�deU��!��Y�km���a�<h�����j{!�G74=t�g���r���"CՔdt!�D�0��P�H�2P�@�#ȝ,Y!�� �����x��Ę�.�j/�$S�"O0��)]��DҥN+.�R"O�Ѹ�-W
��\@N�h|":"O�i�SfE2��q���Vs&!kC"O.���ѧv �)��Y�
�"Ol(�Q��)3�FU�"͕ N�)��"O�=iS�PN=
@��lW�GE es@"O�l��ˋ
�����!4QӴ"O����"զGk��i���p����w"O�h0CjH�I�Z�m�r�;�"OR�� �5W�n`�qmݯT뢌��^���ɡ8����çF�nr�I�cZ2R��B�	�s
�9y��9n��E`�`L�a}�B�Ƀ5d��B��*2��98wI��C�l�d�`�
	(6}r(ū��%�B䉲��iV���9X�تriM����)?��	ԓ�<��3�%�Dq$	v�<����e���F�&l�n�<Q *��`̢Dad�ie�L;'͚j�<�j�K�X��E�N!�`�f�<I��#r�n��D��E��x��QK�<)�d�������b::��y%.FH�<y�E�bUyQ��=�^��1C{�<)�nZ6��Ӂ)k���~�'�ax2�2A�	����I]
U�!�@��y��L�M�I)�%��:l�����y�C-^h�2�,��E�%d	;�yb/V�+���cc�qm|�B�AF��y����'��:��t��HK�8�y�~���q-��]��ؘ���?	�'KV�IDmUu^T�A?�:!i���x✓q���EdITc�r!�F��y��ݦJyp �c��P@N�Kq[?�y��J�4�4M�.x;���,�y"�R%�F�)p�C|q�9��J��y�f�2d���rHH�m�L,�w�8�y���n�>��č��:4�����S
�y��I�.�؉�b+Ѳ0�!�3�S4�?����?1��RD�Em�W�t$�5D�`�b�1\3YҖ臕0� ���2D�	@��gR=2wJ˞=��kW�>D���+�g%���T�Ʊ?D���<D��Q�E�����G�C0��j.D��j�`d�Ey�Bő���o+D�ԩ��]'��<i�D�w�,9�Ƴ<�*Ov���G�9���z@��SZ�QP(_�2�!�d�)d��p�C_��]�'C5H�!�8BbѹI�aaCH�0$}�"Oܥ*�∍>͞�1i�Ie6)�"Ox��'��/���H�RL��"OV̐DI��t�a��J�9t���"O@���tb�1)��'kLQ�E"O|��d.B�8j��  E�f� i�"O�D3�G�{�
,��A؟8 �g"OJ܀�N�1�T�w ���4"Or�I�gҤ@(,����ا8�p蒇"O�0��	X7Kk��T%��E�)p�"O�-+��n'�q���=�p�J2"O*�Y'ʌ�($d�*"��lÐ`d��|�OP!�ƌ�f��T(Q�Xh>u��'���c�陛�.qҔiC�#�℁
�'�����>V>��BR.�"���'%���Q����-��Y[���
�'a���cf՝X�`=b��ϻRq����� hXC�F�^�P)��CR���MP�"Oh��"�A�3�u�@�ۃ�b�!e��ݟ4���O��L��Ί&.St�`	��y.��S�'�ʍI�E�6Q�5��4u�" ��'@R���M��@�u�Z�( ��'�F�P���/(�����HLR��	�'?Б�3��qz�#�ˏ%H���	�'5� '�7��8
���ϖ�R�'R���O�'ujb
��t��sϓ�O����O�1f�L�U�7{��� "OF 8F"ܺ@����K�L��B"O�X���Q5{��r�e�}��9��"OHX�t'��F3��a�B/+�n�I""O�8�/R�l�n�p�mљh��!"OB����B�'���z�lN�U�|���"Oغ���7Ly���U�>�j���"O��b��h��U�lS;D�:	�d"OP��G��+) ����y����"O̥��)̺.��DJ���%6�Q
2"O $I$�N�G	�ipSJ��8���"Ol<b%E7_>>��ɇ�S�~)+�"ỎY���P�F�Z3�M6�����"O4��О$p�i:�M�$�b�:�"O@8!a�ˌea�pp��,�	�G"O:m)6��:ja��a`��%""O2Ԣ��.=T��T'[8�x3�"OF��f�?]F��;�FV'�� 5"O*�q�7q:��s��TD}0�"O�(O�����e[%\V~ �*O���1%E9lo$�pa���"	�	�'�<E)P,U`��5����|:<��'��m˔'H�$	�XP��B�0��'��0N^:P���P�i̖,��!��'^Ԅ� ���g�x�b�g�,.XY	�'�4	��.+F@q0gɋ=��Ũ�'-����AЕ]�ā��+�h)�'~�i�gÂY�v�@�Y�[��,`�'w0��!C�6�4c �)W�*��'@�aP%�9���,Ҁw���'k4k$�ah��KR��.'��		�'MF���=��ɲ�	ʅ��i
�'��\0��݉P&�!ǝ���	�'�Na*�i�A/�e@���ˮ��	�'^e�@�W� �xv!���h�'�0�Ie��h$LP�5o�:�9z�' 0|jr�^b
�Š	44@���
�'�T�[q)H�U�=�p��=a4�
�'8,m�kǿZ��E�d��j���(�'V||�`����a$��3� �3�'=�� cX�A>lBǁI�'P��'�p(Y�Đ�^BJ�q�h�!EZ%8�'E�Y�C��2�8)h�nZ;I�D��'�(��e�DuHi�`�s>��'���CB�ڣR�
&��(�
�'��:rgаCq����.�(-.�	�'���2����H+8U�֩�?d�PiQ�'uLI�2m�-r�lT+.��h�J�'��J�� �"߼H9��_'p���'T,��P�P���I�C�4f�S�'��<W�L=q�Mq7�X�o��
�''|�~����C�����'�"8� ϒ�P�C�f�}���
�'��� gN�-#�LٸUȕu2��	�'����VeJ�-�Œ@��@������� ��wOT�_\���V$�X�"O�=���� 2��y`�nI%s9�5:"Ol��a�7h��gM� NM:A"O��`�\�IN���%�%'��"OV9��AѰ4o*ݱ3&�u	4P"O���
�:�p���[�>%!r"O����Y>2�>�k@��=��Բs"O�  ���0W��зR�F�p��C"O����E�~�B�hĨ*4����"O��J�D�5V,��2G 4 )��3�"O�ڂ�G �	���I7�C�"Or4a���6E���0M�0гV"O�\�f�p2�1C��fk��"O��#2K!4e����7bX&��""Ozd��d�e<���7C򕺥"O�)�7��m��aQ�G-R'
X�E"O<�TJ�6�,	��G&�9��"O`)J�a�7-�xHX���x12�:�"O�\�@�4@��%E��9�x�"O13�_�r|aRa�J����"O�HGfWc�D���@�]�"O�c�d���]�!`@�0�)(�"O3�L�F�������F�0��e"O 9'��,.us� �#�ѡ�"O���Y�M3�	�Q$q�f"O��	�L��P� �#Y37��G"Ot�p���n^�@Ƣ_�P���"O���#��2�\P@@��9�8��"O:�����9�us��F�h�c"Op��AmI/��H*�\<s��Pc"O�y�g�
(��P��1�t��"Ot�B�n�&3�!)��Ԫ°�"O���KͰE����D��bؑU"O4���J 5��#C�%C�<���"OZU�K��b�ؐ��ڪ��0�s"O�0 dZV���kҠ#Ƕ���"O��k��۪�"e�U)��B��	r"OyK3�ɑWwV��2��I�@<�d"O�\�투p�ktMB� ⮵{a"O�0ːA����,��\�LI��"O, �+��x*w��
ӎp"O��dU&B0���!NrĆ�	c"O���L�B���y��	9��!�E"OrqQ�OĊz=���;�:��"O����� "�2 ��@!U~^��"OX�kWÁ�*umꤩR3ZĎ<��"O�5	���0�@U���S�6{5"O��{ML�o[�X�H��:��W"O���J�;B�����֔i�v5��"OdHAoZ�{���3�ҽ}c ���"O�(En�3`e�g٭ob����"O�TpoX�S��Ę3�\�F�)��"O��je�$2ͬP�_�9�b"O��X��E�� �BA�!&��җ"O,yg�	�%�a�  P]���S�"O�p���_�>�(l�礚�e��� S"O����.�2*̪<C��CO�����"O��f(��/落:�O7�@�["O���l4��5Jt&J��N�9C"O�ԙ4+L�j$8����(:�6H�r"OĸƥK�d�j��Jz�,�xq"O�D ��@��1��'p�XDh�"O��f��/<T�݋��Dl$��c�"O�EЄ�H��9Y5��9(`)�""O� n5k�׫|*�Q��ۉ}�L�"O����Y.'��Y󱦘/2�d�a"O��x�DR�=�ĸQE?�r]��"OHh" Ȃ�;��D՝M���""Oް���ܘR}��7�]�T�4���"O~��AađJ)�a� J:���
�"O4�C ���o�rPƉ�L�L��"O��mC51��	
�`�`�� "O2誆
]����q	֘O�d=��"O��)�Kȵ�fA�Э��0R��c�"Or��Ս߻Mx�(�L��9gx��"O2m�09�a�,,jE2u8"Ojsi�>�j�p& �����3"O��q��nc�h�]�'��aK�"O�t�q >L��X�e��|�>�g"O�}��a0Ft4�b���hb"O�����6oz`́�ޔJ �q"OJu	R�&U �S4iYv�! "O&�6B� *a���Ԧ_��"OzL�0O�޼�97�ʩgX` P�"O��˥�/��U�3b�H��"O�`x��j�|�B TT>KF"O�\Aağz��1��^�o���2"O���֥K�[�H)qd�W� �`�z�"O�U0#��|����R��(��ժ4"OxT���O�DRR�[3#�7}zHYz�"OD�;�@"^�`�p�S#5I	�"O��Ì�ji�`���p$dyF"Ol�#B��6��uǕ&;k%"O"���C�r9,i"2&�q�	�"O�)�����k��p�e$�$=7��I&*O����Αn�4<�$G�"� �)�'I^��%�	�~jv��.��C!�X	�'��]ф�i�VD���׾���
�'R��[s�K�{�z۰"��7c.�k�'@��S-D�~��)�pLE�0>�x��'�8�� b��s$�7KM�:ަ@(�'Ĭ@6�����I&K֌ {��'=��`�(_<Woz�!!�1s����'FH[)��lT1gϩir��!	�'��ҁ�H%<�v�"����d@����'ސ4�Ї\��,`*0(ۼrf��a�'� 0���ҡ1X9b��18�0�� ��xҀ�͠�|b�M�..V���%��@Z�o�:txQ��%L2:~~�����	�_.>��)b�O&"��9�ȓLx�h�BAV85���e�@�h:�%�ȓr�r��4&�7�"Ug�G;�hD�ȓ/52`)���1,�՚���f��H�ȓm��`5E�l��� n�6Q:L�ȓR�`�Z���
-�|rb�[�8!���D!��_�**����syZՇȓ�4	�&LL�.4��Z��-�ȓ��[Ō��3~&�6-O�`���ȓJ�D��ˈ�%��$�#�I�cML��ȓK�n��1�@Gl�I�� �(��0��K�����œ�⭳��U�~E挄�EIVq��C�*<@��ږ	Ŧ��	����Aa�5u����7�I-"d��ȓt����͑=��1�JK>p&*���r;2�c�%!�my��T68�t��ȓgO�0�K�`-��3��3��ȓ]t�J�LOR�!#4 P9�0h�ȓs�ؘ �H�,��+�*	64j�-��S�? �L� "R�f�2���(�#�P�5"O��3��B-��!��F�$|�L2g"O�p�R��>1B<�����|Q�V"ON��Yk��Ð�;eB���"Oظ!4ǆG�R�Y�`� &\t��R"O�)k�l��|�A��DJq�X��"OR��BfƟO.���c�y]r=I�*O�e��Ӹi+�K�L*,�"<�	�'�J�+#�/�A�!�89H��	�' 
�x�C�+m��0�Cb���q	�'�8���T�ĩ�DE4d��'�^���jߴXż�2�9� ���'�^���ɵr���@�%�5)�6���'G�ekQe��I����pl� )aHD��'T @���`�D b��\�5Q�� �'$z���S�RT��Z��\yP��'l���(�u��CLŽRaR�{�'�1�6*��u��AS��GU�L��'W���D�اe֘�����l�h��'�h����E�X���f�U>{�q��'�����cЁY6�jvFU D����'��z�[
p�JO�;<t��'3�x���Z FR��y���3�L��'g�t&�$�h}X���0����':��@���h��,r2!Z0!~$q�'b �#m�"s���)�'�3��S�f�6#G���Nq��'����1�Q9h�R�HN
���a�'qrHk#��J�M"a�ɲsI���'����·>	�@�0�:��8��'���cu�-�X5!c�Ŷj��K
�'�}P���2�` *�w�P
�'b���$K	0�Ru�g������!	�'��@p�6fE����
� X0(#�'��,�u��/c�=�LGv��q�'���a�@��sfpA�bÓu�FQ�'z�4sU>n���C�Co�i{�'S�E���^�]�`��c,����'�����g��7-�,�����''@�����%�4! ��p.X�9�'O�����6$!b�B�d�ѻ�'������B4e&,ё�����T[
�'�Q���P�� Ap��O7F9��'�б{�E%1ۚ@k�h�D����'���n�,ظ��w���{~�i�'&ʸh�>~i,l�DI>q��E�'�(���5pAƬ�C�HRN�И�'��kwB8LL�B̘$9$p(H
�'�"�RS�ٹ&��"��6Y���'徥B�*+�V`aF�'�`���'b��Z��A1��\���Џ$���'�d)���_'&1�����1q#H9k	�'�t`I7�� b��`*DgE0U ���'B�p�N�~�I�FJ1ҨH��'�p+D`�GiJ�@��ݜiK�x:�'���JÉ�m,�{dJK�3���z�'�����e���+�T��'��3�ÜN<�M��G��$2�i"	�'�i�%T� {Tu�Sň0�$��'H�� S�U�:�Llڂ�X�$G�Tc�'� �Z"�@�C:����@<"�be!�'�DQ�&ɓ1B�ԐTHվ�v�
�'�2%�FM1T(��jJ"X�(�J�'��bv��M��HҦN&%����
��� \je韒P�0��6�=Bp���"O �
����I�t�]�Êh�"O�4��`خ��c�ۯ(���35"O�T$�Ξh�tX��]�d��9�"O���� �B������e�D�I�"O�1(�A�8
�dE�"n>m2�"OJ�i� ��<tR��E�%t0r`"O@t@���-H�K� �����i�"O�M�E��X��T�L�X��"O@����U�  � ����r:��"OҹJ���)gN�`zS ��K����"Ot���MƉ|¨��Х��2E�
F"O��I�&�'o���"��[*z:9K�"O�DP��S(7J*X`E.��$����"O^a�`��6���mˠl�
Pc�"OxJBo�s�^����w�PtS"OrmJ�$
oZ���J��<�x"O���g�4ʴ��Q����"O���!M�>u����h "^�k"O�(�fg�OGf-[&"�\Z�$�2"O�Xa��]�Kp3�пIo
1�"O�����a�q���O=\P`�"O��iw�;H@�٢x�8YV5��k�̄pC�@2�~h�P�w�}�ȓQ�D(@ԣ����ȍx��E��U ���%b�]r qJ�*�5#-�U��i���v �-?]��4�8<\�	�ȓ$}h�It'�E�$yV�
JNd��ᔌ� 돞	��BboB6aֲ�)	�'Gؼ`��!/B2tC�	�3B�\ī�'p�h�����{���1��aъ}��)�IK?Xú���e\��E0F�AfC!��S�?���
��_{ii��@)���E{���%�UOƉo������.S��8�"O :�'۬����M�+��+��iFў"~n=wvʉ���!J��u1�#ߗ:ΎC䉕R�h!�7�BF���2#\�7�O�#>�yB�;��	,�YP>�%��y������g�͋P�8��+ȋ�Py�E�S����.ɈJ��"f�k�<���C&xZ��J��=�
���$��������S� 8LS���t�8�!��@��І�~�鰢@�<�!�3�K�+K�m�v?1�'�Z$�G+�3k4�q "QQ|�@�d8��<!�O	���IF �K_Z���b�S��x�'.���mB`ӂXq��ʘ`udI��}"�)�	 � �6��̃�28ܵ��K�"�����-&_���3NђH�z@�BmY$��C�ɫK8�@�D!Ǡ �F\Y��5)� B�I��@@ʕd���:���N�W���D*��Rsj�)>*���`���1�$	0D���׀qJ:P����0X�P/D�D@��\�`���u�֫2�ʈ���(D��!4�Ə��1�UH�$S�����(�d`F�<�O|N1r6)��O�Ȁ�&�n�r�)
�'*(٤嘛�d��C�2l̰!�'aqOʑ�ᓉz��:�ğ>i��"�J�9���Is���N�s:ތ냀��-WjX�Ѥw�,)�wn �Ix�'1���"O�(��H
'��=s�� ^ %��La���A�BpQ��#��O��)�W���KZ���F	��C�}R�)�IɍZ�����?�MӇ �.I�E{���'*tE�1-�%^�u/"��}P
�'͚A	�&_��+��=��[	��� 4����ڙ �>�A��,U��j�"O0���Y4g�h��"�[��Q�1"O~���K�*H��U�r�X��4��1��������I_�)�W�8��KT�5���JC�I-P\+�.ذU'�j�� �5���	\؟�R�]�h"-+7i=X��C��.ړ��'��g�8�GϭK���y�i��-B�\�ȓ9�$}�w�W�a�r���(�5d�,�Ih?1+OJ�)�oXT�U�+]ӌ��BX9P )	��O`�y4�E��������G�F)I���+lO^�a��6����fD
&N�N���"O���`d��l���@�F3\����O����	�^
���$�O6	��!C�	>��}���8����,hF!�Eʋ	w�l��@3D�(����q��h�'��>��<�A1D�<�@�	�0���ܧEm� �-D���!O-Ĳ�;!�G�ୱֈ.�IZ��(�0m߀�R� �ꊖ)<��,$�����M:�9R	�D詪g�y���*lļ,�B];j����B
���'�ў�`�Yaj�gڌY*@m��z���6"O�+�g݋up]���+q}�4�	Z�O�*i�u��"ǂ�P�%�?�j,z�'�f�IJS��� 	����h	4B7D��A#L֩R�AZI���S�&5D�`�C��8p��
����n�����4D� �"�I�9�̱����0�K3D����`R -���R	  �Z��2D���j�"FL�\v��>JrT��Q�%D�P�V�,�R�H�N� [���@8D�H�DG�W@0���HP14�(�!I6�	f�����C�f�~�B%O�5�Z\���3�O����4G9��B��Z/]l��b�%U�2S~Մ�6E��n
,�B�Jh
Q��F~�.Rk�O�8��,׎yl!#5��.�q��(]˓�l�'�~���1���E(���#z�Qs�߂E�5��@��bdVH��J�$�� h���Ƥ��$�r�ȓR[<tr¯!+<X���%LjTh8���p��I'��@���w d=�ȓla���MW5�R� ��� 2����ȓU�d���K(Q%�t�E%�n �ȓ1&T�p���R��J��,y�x�ȓ:p���F�]=R�V����@�����N�D<a� Ì;n�ӅBL�����B2x���$a�m�A��=���I\~�	9��u��g�>�	a�V��y�+˺Y�4HK��Y'2M�Х���y��ʳXrf�	�#ɳB+�Q�����y"*n�1Jr윿f���a�yr���54h��&�8Z^f �P�� ��<�U�x��Z�3�OT.L�ڰ���ԅ<ڰ��9���3��6�֍�𬍭-�m�O��#��(ҧEj��E��4r��:a�D�H��A�ȓb�0�3V�[1P��a(�#)Lf��O�OX���A������[$'��T�ċ]q�<)a(�	g�N ���X�N�n̓/�d���|Bĝ�I�NM��L�4Kذ�Iԫ�ynRA <��䌃�o�����A0��d=�Or�C���L �$8�M����|aP�'i剣gޠ��FL�p(,���CS�P�*!��'�ꔢ��I�"��E�/������(O�yA��k�,�a6ʖ�s
�|q�"O��0��d4iS��X�d���j7"O� �$Rf	�1!������'�b��"O�rV�̺[ ��+D�Z9(�,D FHH<�`����YZÈ0} P�]V��0�>���,�d0�O�(U�Ib�C�P�<� gI.Y�*HX��S�o_¡�V��O�<�&`�
s�tr �IL�p�"c�<� #ŁI��l�#�@��$�%������S��yR�T/x7�� W�I]�upRmT1�y2J��|�a�-�,Pfn�8����'�{�	���c��V.Y�����I�y�ˊ�O7z�Z��=W	&�����y�V�4�:t�I�&2�h����y"�E�;��Uڔ"�1"� ����y�M@,|�V�J�����<cGK��HO"���X��a+��_/˺� �.�� !��L4��`2q�҉
�j52l�E�6
O|�h W�E���شi��v���"O�+�,�!t^̉�go�>+0�a�"O��P�aԣ#�pab���'�!���0xm��2P �N+Լ�A��)�!�V�=^��� �^a�j�i1O
�=�|¶��t�(��B'���@���y�<I���\s�8��.��;2e�����<�O>9�Yz`�Sb�A%-���r�� 
��Ʌȓt���M�CbT�3�&�J �ȓ~d�$��䂐�d��sH;\S.��ȓkI��Cң� `p ���I]�}�ȓn.� rkV�a����rZ���6~09���M��x�i����F�E�	~�i����,�ȓNBD������XkS���ȓ!�LicLG�tl�0�C�݆�1�<]�P��!9�Q�J�<�z�ȓF�0��lֵ3O1���愨��P*����g<!���4&�9�ȓ]��x#�N�51�(�VA�5��<�ȓ/��i3퇡bW�!ɑ��>�d-���؀ȡ#0v�̉�5�̅"ḋȓ7X���D�@e�=�'
��Po4T�������+cyr�y2aп4q�h��2���f+^�z`��G�߃s����ȓ#�}�b�(G���w)�|}��AA�����	|��\��$���!�ȓZq$���OC����
�/�X<�؅ȓF�2�+4T0J�N�
��Ώ!�Bu�ȓUֽ���%� qʂ*�n1��7����e������*ńO�4�ȓ@-R0��RMڂ�����7z<�ȓ I�T�RE[ m=�2u� �8��ȓ1N���H@�m�p� C�f�����r>�ap��P�R��5n�:0��=�ȓ>�b5*4�K%s6��0U�_���V�2�`��H'
���PR�n�vĄ�}7�t��Df�&���µD�D��)���a1�~s���Ё�5��e�ȓn�rmIt�Z+u�<˖A�6U�!��FI�<�a��-��Cw�E4H�`�d �����L �sDx��I��2��eT"j�1 B��1WtC��������ЎA됡qT�հ�2C䉑Y���A!� ɺU��DpC䉼D�4Jwa��{|��*g`�B�I�2�<9��S�0����>{W�B�I�q��|�Cf�.�Qe��7lB�	6"�Z��G؄�M���B�)� &xȦ�%C};���	wlHt"O���r���5a�!R$b���"O�`a�%M�-�������8_sM�"Oءr�O�{(�[$o�qyZ\�"O,d�s(�)V���S�*x��"O�x
�띥=@@�m]�&&����"O�$��
�$zt��U��>F��"Ox���?N��(�1��f��#"O������A��K"��1`J��D"OZ�%�۶��mr" ή$��3�"OV���I�>���0�oQ5$M<�1"OZ�� J�G�hD�f.�<-#��r"O�e�#��*��z3�"
����W"O��X�O�C� �XF���,��Y�"OF�`L�;ze2Q����$�4)��"O�q��]|]���6�̇'��9��"O��FG��lD�y6dP��"�"O���S �9  ��QRB�,�2x�#"O,]���?9���"@>c�f1s6"O����*$��tS6Kf���#%BX�<��,O?N������0>���w�FX�<�6)	��4�W��N�.���U�<a�gV�h>�97%��fFM��'S�<!�`M�5[�U��BX5JP��hL�<��jͬJ��\��$�)�2 { K�<IBh�)z�Xx��hљ����S�RG�<A-�''6�BApJ��3%�k�<1Aǂ�)�,3�l�,�\]Z��Tn�<Ƀ���r%	�Ld��E0RHi�<9! ԟGd�;mN"�>�;V��d�<�C���./�h	�#Ή_x!Ha�<ёύ=]$:4 $��ڐ���+�b�<G�� K�r!B�U�8Mn,��� _�<��.�:F�ulL:l[8���"�n�<�vϜ�j<c�D�wiD`R��EL�<A���#����K�-�X����O�<!��W�8�Uh6M���P'J�<��֫+�|��A��/2L\ɷ��K�<Q��8�2D��-�%j�%1�nJ�<���H�L�l�� ��PI�#@�<	'�M�Y����!�{(
%᳉��<�ՂCB�:ę�W���ȣ�Pn��1a蘋=(��抹rQ�L"V��И�� r���W�iZ���4Z<�� Fl� CR�>�㯈V�V���I9ڧbK�%����>/��9bGP�R�(̅�B�p�H�n�y���pA��d���FD��_� a�<�bQ�2��x8�ޕ$hJ�Haa�^�<����3{8�̣VQ�~��$p��8�%�'�O>o ��g�'��s��mQ�Aa$�بx'��jדhU!Z���
0�����47� ��D%@(0�>1��D�Y����Y���b(Y~�����8mڭ�<��	9hĝ�P�O�3(�>r#Ć3����L�)m�2T&.D��
���B�cǋ��"zΠ;4�M�urQ�!��8�~bF��;hF�؋���:k�N_�.w�13GÌ-g�1bKm���,a�Z��w-D6�jP�D�9���2��z�RLslX`D��S��-b�N��m%�|��t*`ױ^)�]�ua	:���I1\.�m��o��d6��Gm�J5Vщ�N6n��!Z�L(h���$�U�Y��L�ƭ�b��H�'b�C�"E
��r,(��O�F ����Iw�z,�G�F���,rԀ�)*���S8�Hz���n��X!��Q��C�ɫm�zP���/rU$����+����V.�'k�n6-J�y5�s�@�0R���$?�S��^�%��u1�Sl�?%�L�k���fh<�2��`8V�0%�K1Y|FA��&wdDaVÄ
W���ݴI�*̂��*�d�h�
Ֆa����d�����<��3��.Cm�h��o><O���!��@j�p��O~�^ԑR�O�a���8����P�'�*2�`	F1�RY����w:�*OƠk��� P�:g��?Q)�ݸ��ٱ?��v��Y�:��&�*�y���z�1��!)J����A62�:dMθ'8��p
����iV���g�%�L4I�E�10h���iɳ,�JIBr�ēE[�'�NA&>��w�S�fX�&��,G���LH�e�P񦄇 �-U��l�L�UX��ҌP�f������lSXEA�,,�	�(��4qV�ܐf��)[-�HU˲��R����V�<�1�*�U����EG��y��=*��Hp��
B�&xp�MH�F͓R��v���@D�A�H����4��6T%,�]�.�D��]� �\�Ѐ�rC�P��c��T�d5sc��23�����-=\�Ea��4L��H�#V���$	h�\�R*S�R�T��p��{]az���(f&Vxh']�/M4`��m�b=��+��:\Ī4��D�#�R�{v�_�A�~���;�m+�nVm����l�G11O����ڜA;n���O��!�hYᖫ��NĲ��OrDؚ�䁜wC���˷Y�h�	�'������:]a �J�X��T�	-o�D����Ӕ$�
��t��
N���r�9�\k�*C�%T��ءr�����"ODs*H�c��qa���8p�ͪ`��5��lk���M'CιX(��"5�$иYR�Z�VvTpF�X3M�ڡ��	+:/��!l٧O����.W�5x�&l���a׭��D!��6oʉZ���y��iC���Y�'�eC�I��]�l'�`S���V�4a����1)vE7{U���w����?��傝w.0�x��ӡ �x$Vذqyƃ	vZ�O��@��hO$� �Q  �$�r1����	w8R�B�����e�b-��D�ole�C���-�B�ɮMRU�UB�<(�Fm��M�Q�	�,�iq�j
�n^n�FD7��~~��!&S ح:0gBh���ȓ�0�i<~�����D�Y"��Q 
 2��(X�OB�|���H���gV�m1Gi�=���X0�.�~�&Kv�i����8�0�` L����]��c�,|�e�����a}"���\��}�PLF)8���#�R�'�~���
�t��c���B=�!��g݉P��� Aa�R���8�n&D���ҌP�(d��[�Pc
n����@B�Z*ʘ�l �u���Ȃ,P�Q>}�Qd�8̊���!U�"x2Q�/D���`f�#+ג�pk�+^U$<(�
a�!��ʙ�T��` �$�L���E�Z%1O$�z�/�>j9."��G�.�5C0�'�%kPIӭB�L���A1�ܲ�aO�b�C�C�<V0�A�H/.�!�'l��ˠ�Y2P�蠵�I4ʠ����)�<0&�G#7p ��A�4�6���o�3.R��{� �i��=i$f�L�=�
�'V C��L���J�h��A�X0y����`bq�b���- LAƅS2��`J�g?��Y��GDN�!����
6�v=��|���AR��e1��'�:�Gh�!���AP�.�2
R]�� هC�O,`��ӵ���'l�k2��W�'3��7�C$��Eb��8 �����c�,V/�����BU�Ș�*<O��6�Y�-����pQ��Q��I�9����r��I{��ܕhr��Co� o�2����PT����ZUq�B�wh<� ��,5͐�V�\,^W�I:�O��<A��c����%ئw�8��p	�-7ϒ�	����B 3m�(�Q�eV��i���y�+�9~����Ě4^�h��瑪H�~�����@iN�i��M;u����~Zc���ʜw����"L:�~hs���*(,a3��K�Qӷ�
.l��'O7
>�toG�0��ْ!�}�,|��{��>�(Oj�!b�		~7���2�\�Kz���I#5���'�K>,F�գ$�9>I��M0�0k ��(�Jh�VaM�h#!�$D*�p5�S`�#dqv)A�*��z �	�-���	U��+@�p�1��� �O�Z���
�'�YR�h����y�C�ϼ�T��"3���+!�_n,2��,ۘC'^7�P}&�����%����]0C%H�S�%���Q�B ɑ��C�	����P!ʦiМ�c,%/�i��
ƬL�1F̫^4B��d�6~�x�(C�Hx��ݠ#�M<!��{BJ?.��C2���P����58���+�	�S�Ĩ��i���D�g.�A��
.ZU0��c e��'T2����`�Z]QF��<�E�	8JN��չS�V�+u��#&�!��M}��	�_�j� ��4EF�2�F�N�,3��<��F1�����D�mq��#�)��t��=�2�U�#!�d�-R��j��O�0e#��O&���"��ѬH�r��T��v}�g�'��|*@!B.�X`��ʻjA���ߓvަ��fIl��6� `r�`��}�z��t�W)^� ��d�O�����R�@B��وD��e��A���(�(�M�"��L�|��Ni1�a��K�Iz�폚^^ ER3"O���D҂Kn�L�Q^rlz�LmI %���x�H-�����kM�?����(��f[����'D���U>��K�:b|��Bc�6m�O� ���F��4e���s2��.��ĂlV����I`��?�(���B\�(oƄQ��r�<���'�*@y#�'���/�kc`�27��a�b�ba�Q�5Z�G{��X����kT'r�`��-�� ��:�g��|���^���Pb���R�V��	b�oӎ���d�?2����s�> �/ʀvT6����+a���!"OA�a�L8�E�$^�����'�r��?��O�#}�Ĭ�Cl����)O�Ҡr���K�|r��>��q����F���J��M�~E��O*�M�N?㟬Ʌ�M�U�x����0r@�$ʓ%N���6%��Ä�xб��Ϧ?Ldo~�����`6�R%C��˘y��kӔĲ��T?�nڸ��C֭Aj܊In��%�(-ʔ�ȓ4ȎP�'d�\�2�h��=�2ݖ'�pEl��ы��4��	�HB7]�n��1���0?QE���|84dȗV�����c+zhȑ"�G�'��>�IL�<H"�k�� (�pMVۆC��>&>@�sB+�%�_O�����x�e֣t�b���mP�`"��I��/�~CNf��h��}i��P��XD��I�!N���"OH9�v��1��Ic��1�>�㣑x�.����X�,+1ǸX�C��,�T�;�f*�O��PߴG'̽e�:�x�ē�pI�0�ȓ;JT01�ɹk�BL��׈2����	s�:��6�|҂A6\X�Y�0�J��	��yR��;�<4��	�x, ��G�+��'��DyJ|�#E�2����wQ7)���۴�Pi�<�ڛbS^��v'��;A�*�e�<qE�%\�.!�W��P��		#��c�<����[�8-��ن�t�Ec�<i��%G 4�z���.K6��gm[���DSY~B�o-�K`Ǖ0_m9s�Հ�y��d��Ԩ3�p��R3��0�(O\ۃ�'�'d���%+E�ܕ�`CS� nB1�ȓU�����5'"r�솃 �Z���5̄��GC�;�:����Ҳ)���ȓ[1(e#4,pA��+D
�2h؄ȓ�p-����u���ˇN6F ����}m<5 ��\.+|(�� �f���#Ӏ!�GNܠG�8i��?�
,��b{�<FKU!\v(5�0g&1�fņ��Y�(�-X
XlCW!"�<��X��dIB�%=���Y��	V�t��ȓ/���B7*H�1梤b咆`�X��m��$���^;J�[�P$��U��s�� ���	{zR%������|�ȓHa6P�2�d�jMiTCև>�p��l3,!C 勺B xI�b��}�`�ȓ&h��˔�^�N��|i`Ȅ�N���n�N-at��Gq����������C3^mٴf��tQ��Z �� p��M�ȓ��#C�L8|��J�l<*�ȓz�Hs��LB�ir� 	$\Ј��O�����&\�u�0�$B��v�|��>��h���%f�@���E�݇�+a*u�F@ܥWi���A�\8�
��ȓ��0�대�dݹqIǂ"݇�^~T.[�V�=�փ]ȪL��S�? ֑q�2]3��[�DN�dA�"O�+U��nB�j�c
I�,��C"O:����BP�y�o
�)Q�"O"��0Q&z8X���x����"Opص"R���)2f& 2�1�"O��*��G v{��yF�R9z�"Oz���Fg�IQM�5RE��"O�4�c��I�� �e�":�Th� "OJ4 ʑ'C���g��6B��H��"O�u�B���O`t��[E�6��"O�FcOY6�HF�?:�<1` "Oh����&<�}{���	4>xC"O�r1l�.���#!�؏.F��#"O> "���%-Z4�Ԇ�93��!"O��%��*Xk���N<�|�q"O:��Ib;��T�*.+$�ف"O ԉcaэ��8�r��L8 ��"O��)�䀢@o������s=t���"O�,ʒFC�W_�uqTa�0���"O����-x�ğvhN�"�"O�ivZp@qBoY7�:��w"OД�bi� hk-M� J
���"O�$�%M�ƙ�S�U!$!zܱ1"OR�9r�[F��	ijW�Q+���"O$|�P��.��< v
]:���[�"O�a��3G�5�DCů�đ�"O�)Q�;F�:��GK�_�\�S"O�p� a�:c�4�ʦ��]|0@ہ"O����%H��$��j�%z�( "Of�Q�숵�v�B��KT�E�"Oݱ!	׬j��9B�'^D>1��"O�4@b!�4<Ź��\�d����"O�2A�?X�Wʙ�)�rHKr"O�é�24�� ��@�j1lZ6"O0mb��ѿpX�H�j�>9$�9""O0�k����}�^��pF�3m&mQ"O\L��O�,l�nL�G˒�2ƬH"O�P ЫĶ*�
���J��f-��"O��F���T�h(*��	����e"O$��oĉUp(d*5%�!G��"O��Eh��#����S��=�@"O��ivm�T��'k�xA"O��b7��+?�j&��7C���"O�HY��R�5
B�N	D!$���"O����MYCr� �����9�"O�=@3�Qv�� ������'#�Z�!).Z���Z���BR�}b��eK�:L!�Ĕ�y�X�pIޒ���c�$��d��O� )��Y�QGZ�ы�)�)D 5ʃ�N;� a# �r�!�D�Dv�jc/A3Z�`����P��p���5�0�'EFF�,Oh�JDiB2v�8���,Fn"D�"O��AQN�
���)С�Wz��W���$h�0-N�b4��	�[���L6KP�1NIooL��čp�3RCZ�Pj7mR�e�|��1�5F]Ը��q�!��P��>!CCǒ�@dl��h�(Y�1On��(��^�U!M�r�O`F��PM�� ��Ek�E'21�e��'g�]˲�0��q�r��: ����޶*�x 8c-��A��~�g��^.fވ��a�A[b�2Q���C�	�
�E)�)���B�8���Vv�� �ЖG�6 ;�/U��a{�EF�O��P4��~T��K^�.<N�����fd�r��-:Du�ٴ?�iV���kB��豉E!=�.�ȓa^D�͐�Phb��ܩ`�R�%��0���*g�L�I�A�4�h�&��T���[W���he�f�@�"Ole�b Q�J��3F^w���c�LW%*
ـTP� B�p�g�� *ʳ�D�l��aB�'u�\��O�]�p��kj��򯏵[`��PTD�$_����X�.���pS���|}��S�����"�)�FP��ϣ&���p�)<ODX;�
"%���P�i����FT^��\���2F,���'?�dC0g�p$����B����9����Ƴ˒�Ʌ�F�Θ��բ��������0u��sA�Zn|�'�N��J��К�� ���g�a��I�4��: p�ĥ�HF��J��'�@'>q `�ƉJ6�&��X���d��Q� k�'6�;Ռ�[J20Xe��pX���3h�"B�X��S�I6X���*4�I�(��@UꇞA�*
՟Bڀi�"\L�4dʵfB Ջ���M��$r�G��yrN�`	��x��G���(@�=r��1RF��%�� X���pG�#!r�����8�x-�">*�t|���
�<�t�"O�i0gI�%L�e��DQ�7(LJe�u��x�T�Z	H9(�çQ\�y �	g�'�����[4o����&��Jh�	ӓ6^�� Sa�r ��@��<~����._<Խ�G	��}�ga[�l�����'����n��!@��a���}2�yBؕ� MbAkZ�?�<�ba┭Q�Y`˱~Z�k� *f�ix�e߃8�i�櫑b�<�t���/� �fEY� 76=�dRH��� "iT�!! �A E��t���yg�Z�2�����$�\�����y����3���s��9
׆h��Z�S��q��?C�4�o�0TT�R*��2o��(��M�N����t.\$a�1Ae.LO�ew�R3�:�'����Ƅ�&����&��J�l���'
��4j?I����LKJ
("L>�,KI<4� ����EP?ˇ'om�q�`�l?a��%�O��Ư36s~��G�S,�ȷ.�:>5R3��)Ѹ'�����Y�,�ηL��xd��0 �Э*�+B�d�TJ E$�b>U3Gխ&�$5�E˒?�X:0�7D��ٴ��+�85R��
���/��И�A�\�r]Pw�>E�$$ƨr9ր��O>8�pm �D��y�NȕI�l5�� ��?]ڍ81`&��5x��{�"�N�ax�ɗ�$�� #˕�\�;@� #�p?1���%Y=R���LK���b���&j1�XJ"��ϰB��f���b�@�s}t�ʕh˖���>qV�/+����O�d�P,��uWE<<���������x�V>�y��Y$�hPB&F&z"n�S�M��~b� 6;&�S�ڦM�g��l	D��i�	
~�	��"\o�4�{F�ǃ�y�/�`�������g�(���Ҍ �и#ƨ�*,H�[�m�+	x*� J?���d	5�r��փ�t�(̱��^�a«՛oP-:�/˚Wŀ��r(͘����"Gӣ2���*��5S�Y!�������
��X�{��
�$��E"��4��*��s%��O��+�	�-U��u��ʟ_�0��V�8�1����y�E X�����a",��9�M׶�(Opy�&��#^������i��$OD��
I�M�N��k/�!�B�Y��ٖf��L2>4�꟫U� ����I�keR���>E��W!@���&4MDܨg)$��ȓp4t� 艖O|��H���S�2��@K�\���G@p��D�7l��q��=x?	��C��@��|2�
"-5"�M�'eAL�B"iX�Ő`�j��ȓX��pq�Ef6����V='��Ez2@M-IvZ�(��ӈ�Ԍ�BS:j�:�+sAY�2�B�	 ����借#Nd���	���ܽLS
�1�{���5��h�w�Y�J�ЙRH��<�B�	�:�PW������L�B�I#Y��h��UB�����r�������{����'�Zm��1N���ۀ�+C"��j	�'�b�
�C� (�l-S�I�E�hB�����Am��R5j'ڧ_|%�B�Q�p�������%nl��l���*� (@
���+�#K~�Ӧ��.a,���>i���O�I�`횁t7VI�D��\�D���"OBQ9��Z?Bz40s(�7��a�2�'�������7��t���G��m;��Z�A�蘃Á	^�B���θ;���uȄ�M3��ɕ��<�����r�A��	_I�<	1e��`�n!��u�X��@`�m��5����K�nĲ#}�,]=-����Y d�� ��e��S�? �{@N��8�v�ɥ� �A(������L��S�G]�D!�g?�Uj�, ���'�z1�e�Px�<��C: 3Pl�Ð�~�Z\������#PD$K:����'l�XaÊ.ZҤ1���Ks�@z	ߓ���D��%n7�&DM͈HH<���)��2!�DϘ4��;&�!ԾТ֩L�$��y3"�3m|mE����9�RtȰA��c�@�B���yrID�AL�#S˚,��`�1��<�F�
�м�����B�~���
��P�1�ykd����yBJ��y�080#c�� ���J��C��yB��.6>�%�e)�74�i#����y��ǵ^�����);<M�b`]��yB�Kw���¯��y��2���y��X^�����~�� ڌ�y""ќn\D���Oĉc��D8�y����~�^!����))'p���y��T�H�N�3w�L-&�$J��#�y"o��Q�X����<k�쀲����y��	%�.��m��)��p��y���� e��(0�� =8��ʗ�X�y�fY�&{��a ���Q	�m$�yr�J�,,� ȵ+_2� 0�f ߇�y�-�8s�䭹u�= ӊ�zF狩�y�bܐQ����5�,xVv��5c��y�IX�I)z�3�L36+�ń�y���AyDܲ4��g��)�y�O��#y@�Z��C�z���w����yg��m�0����Ly�(����'�yBD*oF	bB�i�.\�`�\/�y���u���dF�R�h@��#�y�P"Vt��f�E;�����⑍�y2��fH�	�_.a�1Ig!�͚2��8�ba%(9Xhḭ̈+J!�ɯz�p02t��
g0Ԁ2�L�S!��0>��C6�>-�0,c'� !�D�?O~�p�AQ t�$�,ۜf�!�D�/k�9�2BX�
��P��]f!��ͥ4�<�w/�*
�d�kÎ��SZ!�DD=~q����B �+��5��Z�W�!�)��E�Ab�-]��}��m��!�$X�f�V�� BZ>L�le w�4�!�I��-ub��J�2�!�D&*gQ�D	Lif���mڱp!�d�7q]� �dH�q�h�)k-Ln!�/a�������JVx���Q�<�s���}����0/B>�PyIg�FQ�<q�S=MN�sAU�q"t����Kj�<���9|0�AV)ɂ>�T��Bi�<�aܟz���b�C�9]d%�e�`�<��H�rz$�^��R�B���^�<q�OS&���a&N»e��b�l�_�<��+C7��MQ�F�K�H�)fNPU�<�0"��,Y{U(΋/��p�d�Y�<��T" ���%JB�.D�CU/�Q�<��#�<���'��,"�U����O�<ӤS�`�FX�{}$��NCm�<�uZ�:�F���O�t��ݘU�R�<��NT�2\ĢQ���"Sg�<�A� 9u@9�D�._xV\0���b�<y�I38����hB� i�٫
�p�<��.p%z䆌�p��\a��G�<���y�`Pxӎ�G�Th�n�A�<UI-�� �'d�X˴�����x�<q��N�� C�_028�S��|�<� Z��lR�{'ҐjWe�0}�>u��D�L�8�����*qZ�0���'�>%� h�??�Bљ�)އI�m[�'s�� d���5�4۱,�:�4��'ʊĈ!�B�g� 5���B3�����'%����>�$�S'L$\n��'/d�ہB�J����p$����s�'M��pn�:��D��~y̨��'��yHT+�zޥCP��j�jّ�'��!��"�f�ThB�!H�N�@�B�'t��(��0 ���p�}���j
�'%�l�@IB<��Y�@ё�PK
�'�>�X7�O�!��mz������B�-���?�$�* c��H�ZIf
��D�r�
"��?{�V�M<E���G \��tp�O��������shz �u/��ēl�a�C�$��"��JQ
ܞFr���1@�	��I8=���;ç;A,|:�^3d=j�&E ����O�1�;5(�th%�6գ�]�e�X��M
�-�n��U�'�aQv��;`ڦ�Ѳ��"~�LخWf�y[���0``�,�@�h���ru��7e�	f�b?E����1�U��<j�Ʊ��G���X���_3[dȫ�M\;I��	���O9�Ѥ���Ԋ�9+d&� A�L�%n~ ��a�H�z��RFB��?Q��G /q���B<Y��S�3�!z#�W2.�j�� �%�<�1C�'�x!��ֻQ
a�M��,Z��,b�ґ0ԡ��H�640�'���*�]�CHM�̟ �?uhs�Ȩ��Y�GיH!�L;Fട�f�"<��@AF���a�hG%8�jp#���Sw�m�B뛼�M�g�nx�g��4����m�\���@[5t=��J�aR.������������+u2�Z�/�:���.i��C�ɱ+��MZb��7!4�t��>!v�C䉅$�f�C�G���F��F˃N^C�	'd�ڥ#�e
�$��Ҵ+��"C䉙+%ujU�2���%S5C�C�ɕW���įZ�t�׬֤8IPB�	O�0`6$��0�P`sSJ�Q�8B�I�;Y���s*��j�0�$9��C�	�:�h�S���</� � �,��C�	�]�v���D�1T����o2�~C�ɮȠ�c����.D�
����=fC�I.���C�I��m%����oFK�C��##�fљ�M;wb��R��9g�C䉪Oj�U��%� ��Y�p�[�1�lC��<1��a��R��� �1�U
�<C䉈K�"0�m�ذ��T�	]�B�I!,ҹj��
1r�컡e'd�fC�ɱjf$�k$l���~\�"(N"C`C䉷!�*�

��H�X�狍BZC��2 �:��W�ۥ"��"
Ǆ�C�ɰO-�R��AT����J^�B�ɂm�@�1ب���a>f��B�	8@V��Q�Ȅ�!����#��(G��B�I>�ز�L[��: �*�5,�B�Ɋ��l�b�	"��B��>"��B��<M��i��`�52����΁cw>C�I�&l��7=���tK�*p�pC�	����v�
�
|��`�X"N� B�IL�0��0k��H9Z��U@ɎP� C�ɏ$z�(*P ��Sv�B�
6'�C�I��X`qc#�6*�jT�U�R�C�I�0����GY�)�h�HS�t�C�	��ܜ 7��������$U�C䉭�����xT��;���k�0C䉜z�87(��Q��t6��C�6J��yR�g����æ$	/�C�;N�=��e��9�lʠ		 �C�I5N�h�3�FJ�P�h�H���B�I&fu@f��X��l�6���5d�B�)� ^lZp/܎@���eG@!l�jm
%"Oz���P骭!P �X �tbe"OPU)��8a�=
Fl��`d"Od�B��m��I���K�y�X��T"OTd���qs�qq�g� �:P�%"O��	1�L�/�1 ��`�.�0"O:x��I�-
���J���=�n���"O�Y;hB�t��x��ER���"O�U���!r��W��� �5"O�`h$�23��|y��:	:0 	c"O�	"�k��e\�����.�H�r"O����0l�XA�·� �.�ɴ"OX�� L�U�&U���J�9�p@�"O�(k�st,{֮��v�8���"OPA���E��L|*f�
M~>�#V"O��v��/��������!�"Oy�$үL�n�H�&یEa[�"O�9�F���"�pQ��~��80"OL�P��Մ_���Y#(Tx��	`"OdE�4�;u�6sV	�2P�\9�"O|��u��@p��" 	��#��)#�"O@���
�Xȶ���y BԂ�"O�1P���Gz�ys.�r�>�)"OR�q��!a��`���X�)*F"O0���NLvDfq�-�n�0"OZ��!�92�<+�,ݷn���"O���P��l�`�����,,ު�J�"O&,�OP7jFē�凶L�,�!"O��B�Jx��A�ʨo����F"O���!�
n���C�� u��"Op�c�G�$.>�[a�^)0�d`�"OV�����<D[�xKa	��^�9X�"O��� g@�&����
5@@�6"O�\�T��5Vil��å��}R�0�"Oh����~z$ ��5����"OX���P�%�����oˠs�6��"O��a&_����m΀`�$X*�"OHX���1`��$sT
�+!p"� E"Od���ܷm\.Ȣ#�9a�vp)�"O>�Q ,4K���p�M���"O�0�F�8+>�L���N+-(���"O�	�D��R���f��x��3"O<���#�
�@hƘh��@��"O4��W	WG^Bp��V�$
#"O��2�U�o��l[w��D����"Oz�j2�˙g�8��ذ]�.I�c"O����6�4T04Ƅ0Հt�E"O�A8b$H�\Ķ5�V7��k2"Oz|AS&V�Pf��eaN�RPsc"OP�k�0��B��)�6"OD0�5N�7��tS�̷\���"O|��qB�� >D�Pژ���s'!D� ��Z�Jܨ����ZP����B?D�4�C��Bz�y�
F�T#�ؘ��(D� ��O��[����BG�vY�00�2D�t
Q��9 r^���Ϙ5I�v�j��.D���2+�H]�{�5����n,D�T�A�
CV�${E�.O��$xc�)D�K �]`6غ��"e��Ȧ�<D�H�t��3(�C�&�60u�MAO%D�,�A�߭[�(�i�4����1)6D�x��ĝ�@�:E'��Ī���3D�����ʦ7$�P�ף'.2Xp#��/D�	U��h�<Z&��
2u\Yq��+D�� ���A�ڀ0��Ǆ���01�"O�Xc� I^�TDHD�׫9-^�*�"O�����0+��B ��j�P�""O�����D�L:3���U�t4�"O��rB��n�؅�r��_�A�u"Oz���
��D����ߔN�0�6"OL!�tɀ�5��ݙ􅜹Y�Ta�F"OȠ�lƚ~���B�m@*�I"OJ�@P�V�(�)�G�,(Y��"O���ġ?=���G�cz�5
"O�,8F� $62��@1��T
�"OA
d��"�r��^Rn�q"O�Az�y���
W��2k�"y�"O��[�J�ST���)7��d8�"O�̘����ܤ�CO�R�X��0"O�$(q.]�CSu�/.�D�"O�qA�&n͖���j��?)$��D"Od��� 7���I�@n�Ĩ4"O�}�0	��08P �f�̄(}�q�p"O����#�m?d�Y6N =n����"O�}Kv.��\!�A�Ӧ/:0ibR"O���LzkB�����# �؝��"Ox���CX�{o<|�b(�[�4$�g"O�HZ$��%��9Ve[�o���"O$	1��'����b#K�?�*�$"O�g�� ]H ��"�)m
�s%"O\����9�*H1�@_�h��"O�ԓ���7oT�uE�JUq�"O��r��ϳIM���@f��&}
94"O�e9�e�$#�`���bmhT�G"Oj�*3��b��a�a%�\�E��"O���я1�p���a�4?a�Kd"O�Q`�)\��RA��@�aCƕ��"O����0Ph�"���>���3�"O�M('�P<&������,6]���"OPa)Ӧ#$5��$�-�]q�'�\,�$�H)����Ká��\!�'gh���
?D:�\Ha��?>�r�'z8-i$�ӿ;+�E+l�3���C�'�6�@!��i���a�q�	�'޸łS�%Q��� a	M[3�H	�'�&Ų��\3�~�X��MO�p��'[&���ńVe�<q6�@�O����'�d�B�gٮ_`F�25ᖖA܄���'�fd;�O�Z����Tj�L>Vl��'p��(vR�%���5$:<��'Lj��AA7cmJMK�g��_!��'׎Y��Փ$��Ū��u����'��Q"g�χ>�Di2�Xݞr�'8�ʢh@5I�zIE��!U)ਨ�'�v�:�Ŋ6*�:��5n�9FNE��'-��as*� ��[f��;��P��'��	{�oH�/�t�����2�l=��'J΅�4�ц����͇{&t%K�'t0����o��`��{wD���E�h�S/���ڸ��a�,@ц�|�24�A�P.�T3X�}�V���4$4�vԞR���IR`�)��0�ȓ7�t�wf�(�uaF)
�i*�C�I�5�^u9Q%[sO����=�jB�	�x��H��5.�HAhO�z��C䉗|�tP�6�l���t��~��B�	9�5yg��$v�K��G�{��B�s�F ��)Y>@=�dŬO�hB�)� �\ap��F�P�ʆ�1���"ON�Q�,ޔbX�q4I�6C�,ț"O�i�6�'|�`nۦR�L+�"O�5 ���*V<��=3L����"O�<`��	�	DD�^�[6.��w"O�\@Ěx��`��c/N���"O��!���l�,�Q P�\h\�t"Oj��cIY	�.��$ �����"O��yT�Q��@|��67fa�%"OH4Z�`�Q"J�
��~/�-@�"O������vz��J��ؔ)��#�"O�p�J�/T�N�2Sń��U"OFx� �$�6�!'Ϟ��ċ�"O\�KW3�N�2��;�����"O^-"$K%G!�X�7����
E"OHE�����>+��;o�o.D��9-�729.(��&:Y�f�zak5D���UK�m]��Z@L��y[�h�F�3D�t�4�L�k�习�㙖7����?D���!	�Z#�]�c�\.EY�2R�<D����_����88 ct�<D�piA�W7`b(�Ěo�r�a�j:D���G�)I4�& ��i��4D�̚����'��=֥M`�@y�'4D��3�J�(و��C�M�i����%/D�L�3EP�B���Qg�G�-)��m+D��÷ K�%.�჊�5c|̱��>D��Á�*%rՑ�B� �f��.(D�ذ&��j���	��_�!P����l$D��z�+���#ə
�ȡ/$D���j    �=XR�|8�,�ٟ���؟Ȃ%�Ρc�*��ÑC+�i�R�KΟ Ap�%?,O�)l��M{R�K?��i)seT���H/U��Q�A��$ܚ�3��U��#a]"+�	B�l�>������I��p� _�\�0p	Qa���T>d����'	2�'�A����v��OB�'��Dׁj��(��%G��҃�8;�V�"��ū�Q�\�Iן� u�-?i�'yV�I�K�`AA )�(�x�B�
L��*��/����Eۍ�ug	S�����6pn��[wyBHVN[8�P��ƭU���Q@~�� �'H�đ(.��2��O,�D�OH�iV	b�d�����=+9L)xm��SJh�¬�<	G��&L�h����?�����M<���R�+� Bϙ�G��A#NA~Ŵ��?��=����#�~�f)jN�]�hR�E�7g�p�a_8]jd���ǣ?���v�Vy(��Oh��C�uy��OAX��:OJ��"��G�8U�-� &��tY!H�OD���O���O�aE���6���?9�d�L��9�"k���[�$��?y��?��+Y~RY�H��ҟ�s��L%+Q��{�Ĉ�=�h�*Ď<32�|�"�܁��0R"�K���'F��+T�n��4hT���'������gU�Mh0B`�7,|~L0�*V�J �!���Iן����n��I&?��	�w���jŘd�m�(O�<O�E�������%Ole�6��ty��'�"� �~R�Ǘ>�h�hY&���ڤg��8�l�j��b��ӟ|�)<& X�;@}���'ɤ������tQ��F�N$��Y�dL�m�B|���n�*OH��ɜ�����ڟX����h��4`ŻGA��@B��47ƽ��'L�U��i�o�\�B8��ן����?I�f�
�dT��!�H�Ȓ#g�0((�'���П(�I�x�d��$IKN����O4�!r�O?Kx$!qN�>���b��)
7�M���"v�Y�r2O��2|����&b#��'7��Zfޭξ�b�蛖���I�Of�(���1�D�O��d�O����<�an*W$���D�/�re0`N�$X�Aq�@����O��$�M���By��x�B�R�P3/����4�ޖ�!��D�1r&��</����4y�ɢZ�Μ�#��(Q�"����dH8D¦J����X���Ms4�'Vj���6�'n�O��3&�?1�u�[a�N�@� ��ػ�!�����k�e�O���O����(3���O"��`ލg̞1�gA,	�Tu��ȦYy�4D���fZf%�C���?-�:i�I�;��"dO�:/nx`�B5B'Vh
$�\+7O���5Bt�ɧ��,
*O���I�D=.����ԟ�&�0H/�I1��Jm�AA�p�Iџ���\y�ɛ�]�y��'w�'٪!ʑ��'졐vjZ7Ow���t�'�D�j�O���?9��Q�b���d��`d
����(��N�;�qڇ!��S��牋mh�tRӇ[�}UB��?-B��O0p�4� a�2�[�l�d�}q��xM����?���%�Nmq'��7��'�?���y
� �t[gS�	�"��P�_
Q�z�:a�'3�����27�	̟��	�'���y2OB�0}�T��J��t�E��C*�5�!�ߖ�?�3LG�.D�[w \Ȓf��OJ�R��V��u7��p�p0C���T�ti�ӏH����b�xy"��O�t�u'&̐�D�O�D��4`؁_�|hnԔl�Z} 
�5/pR�rؠ(s��7�?A��?y���2}@,O��{F�A�x�,}B�b�buH�Quʵ<����?g|?	 j۱k ��'+��}��%���ɻ��@�0�؄ˀ���F]��CN�<ょi0�$�5�e�<	��'�B�c��ݸSL|��e�ЬYv�� ��J�	k-"6�'�2�'���'^�	�E����5��ޟl�6şS5\e���+T�b��ujޟd��ğ���2?*O�IlZ��M��헆!w��Ԫ2x���I����.�Fd!F�Ŋ3A�����Ȝ�?q#g]�;t��]h���0O�֝)�y�`�"5ڽ���8p�{��B�k���	#|����?�����Q�A,��'�?	���e���*�+!�x�F���?A���?9@ʚ�[M� ����?����?��^O?1�
݁ju�Yx���<��<Q�ˏsKl��0H��������X譯�`� y(�'9�A�A͉q ugd�ڝ�I>I�Ҹ�I!6>6� .O�h�	2aJz���b�����I㟌 6Fןk]��J2pn�gDJܟ��	Oy"�W�t�~����'=Z�MC��cg�u@�ŗ�K�ֈzG�S\�͡vѹ��<�W�i��6��6��$L/�`={�Oi��ݕ!��a��a`�X��a-P�>lx��w\*4ϓ�u'���?�V��>��I�1|A!#oO*����eJ���8��pp@�D��?����?a��?/O�U��K!&\hc��+t&�������F���c�<��?��^~~���`�	�-q�uc��Jy訉���O�\��Io�$n�x0�ӊ6�t���lV�d���@/���D���J�'�|��@g�)�����'' T���i����O�wxY ���O��d�ON�	�)�4�',��jB�Űl~����K�>)����B�.�I���?e��O1����y@�xz���]��D'�߹x�F/o�@��G�O<E8��7E�4�Ov�Tnڜ~
~9�����?p%�b�-f�@y�l�? ����NY��*�-���!S����8�ʉ/���?Yo�t��A��;i�ܗ�s� i��ޟ|��䟠�'=t�H m�-*���'��!v���k�cN	w�}be�;��ަ����<�q�i��6��!g���ش]�>@Ӆ-W�i*�r��۠#�l���7v�"B�g�*�ꀇ[�����'&�.#����u5^�#���Z��Q�K��^@{Ԋ����	ݟ;�`�}Ő�'?y�I��u�&�:W���i� �*ze���T�z �0��ޟ�����ɥD���y�R�b�� Ƹ0jh� �e� ]�V�:����>��&�d�"��$r���1�'nC�I�׺ː<���ۀA��3(Z�QF��X�J�<���'�ΕVjѻ�B�'z2�O��x`��Ż^�4��@��CT<�l�h��i�d�[]����O����7�����&|��A6L~,���Z�y^���?yڴo�(��H �E�w-��?���:kJ�4���� �MI�� 3J�T��#D�:2\��e�~�,�󉊙8N��(Q�˓Uc�ϙ�}������<ϪaY��$"P��a�����'���'MbX��27D &��8�	�Q�X���P;��sN�
�L��	П���	������KĦ�ش����-�#�P�#F�����E�ԽE����D�0+��y;z�[��w�-Y�L̕X�~�!��w�u�E�n�d�Y�@��l����,^rha@���?i���Bu�䧕?�U%�f�FL�C�ͳ8��a�lI��?y��?�Q��+�9p���?��?�f`?IVLӂ`�2d+�g�.(�� �uH e��I3a@B�� -��-�Sid�p#�ǂ3EP��Ƀ�6U�w��]�\�W�Q�Kl���S�I9{;R�%>~$˓X����7� ���'��'<�T2p�%���V@A-�x%r�'��\���"zZ�����$�I�?�G�<)SRɂgPbЂ,��h#�\��'�	˟ ��-x(����#Pn,�ݟR�h�d��|+��z���qz%� ꘞFF�"�b����Q�'��NNQ��K����I#�U1Cf@"M�HŰ�� w�J���~�JYx$��/�?����?9��?-O���N�(w�T�Q�$_'1\9)3�L��h�	��<���?�b�JK~"Z�p�	�8��;F�Z�~1Xpb���?nD����c�,�s"#�&��Dz��֟�+3�R+~4�C<Cz$��'�X�ȑ���h��_0�MzӾi���$\�5� =*0��O����O@��P��'gN�@��V<vK�,Z~��U��z�J�l�OH���O��i�'���?Y�w�"|8t�X�"q�ݙ<�a����?����T?9tgԸޠ�I�?���J���٢���!�X䡄A� W>l��	|���ɞ-H�\�!�'"����&�<e�'��U�E�Bv!���r�ڥp�	A0��	�����'���'��ɪQ\v�P�O���	����d�ߜ
(�H��&���i��\�TSd*>?*Oj�D�Oh���O��;B�X�(=��B	W	_�5���5Z��� �'֬���/�8R�uK�׬�yB��ڭC��'����Ҹi�f���KU!���E?J0 !���?���iPx��k����'�?����yBČ ~}��tҰf�u`�D	�?�5c�'5��tx.O��d�Oz�3Q����dKL�A�E o����AG�M2�0;4�ɭ;!���ɷ _�@"V���dK�14�Q蟈K�OM7�Y�Y�` i�b���n=�'.3k��:R
�+����� ��/	)�>5������?���Q�M�	���F5�A��'F_����'󆩲��L$N��'��OvL���T���u" .���Sb@.n��!g��sy��nӲyo�s���	�:MH�R�L�x��I�C�<��пl h�se?|"�D��-�;�ʄ��7O�`�K�?C�̳\剈�?Q�/��2���Q�!��N�T�R�Ֆ��Y鄧�?����?9���?a,O|��0������Q�B����`�yi��@��+Ʈ�D�OF����Rq�	zyR�'-2�K��h�2Ď:�"����9SC�Y��I��#O�}����y���	^j���fU}q�e�|b�4�Di�Z�6��s��{+�y��*5�T���'��'~�d�4k��O3� ��!���I���7��6t��Xj��'mb�'L2��MO�	��	h��I24�"c�k�`���)+"�4a��O�S�
sG��O�6��-�5I�����'M�ј���8<؉D�I��q�1�Θ�	��Lx�/O�i�Ix��Q����韸�	����mWGA�H9P�O�'�:Ah�%����Fyre��O �}!Q�'��'����9GB��y�d�'ԡm���3rZ�t�'�r�'��!c�'u����K?�?yW�S�*NfHrb_/!|H%��k��zA�UI�-�5 W�}jt��<�_w�xi#�|P%]�T��b��r�"E����f����@�R�?9�]��9;���?���?�����T�yi�	�gAX�\_ε�t+V/F��a�/L�h�˓�?�j�2 �'��	ퟀJ�cO�e/�`  ��4/�������Y���jq���&c����ɀ�`1(P���:��5�y��p�D��g�6>Ґb�&�js����O�9rs�Co�����OF���rH��$**#;uc OK�6 �ݣ�)*�s�����\������>>�u�'�7���,+� ���_JR^	���'1�
��~�H=,�+��r7J�<!�@9�W�(#R�z%&A,1�<��W�}�\���VԲ8��h�OT=���SPy��O�!�5�C�p%~��-Ψ��Ď�ФY{wNK�5����On�d�O6ʓ$~ի'ۇ���O�0q��U�\P�)�Aщeo�l�e�O4:v����'z��'�N���'��ē�O	�S)���b��#4 ��WB_�]�>����7(=�ӄ��w$��"T���;8n���>0Zb�)Ɛ	����bO
9��2R-��F���'���S�"�������'��>Ot�&��OJ� �!3ㆉ���'-�ܻb��S��ן����Gؖ�y�ŕ07���A�L�V(|��Fj�7Ъ�Br���?���\�OP����L�9���U�n�QV�x�y!���(_�<�#bÔ=/a`MK�$Y�P��PE]�x��� ܤyĦڪ�?Y��?!�'P�,���\	0j��S�NRW?>�Pb.���ѩx|�����O����O����|��=�.L��̎�<,�ź��8:+Or���O\T�a�O�0���9���E�nh�[��:{�]s���4N
,�t�˼p�<p�?O�����?YW�C�,剓�?��_/`Hb��W�C�>Չ�/��3_�-��θ�?Y��?Y���?)O2�������d;%~=r��P�h��'�A�n�$�O�d����ly��'�2��*q�< pfM:H�*y�D@�,�i ��s����܇�yr��BF(��E,v�P�|�35���KvH�4�bX;���*�~�Ɇ���6��O��d�OH�	�ވ�����P� X���n]�d̬���
�4����O��dO���2�<����?Y�D�c?��HL�� ����T-0���:6��I+E���7��O��	L�4h�\{�$#/�ˮnbj���ͱ��љ�ˌ0)��y��m��?���<(�'%N����� -�O���O��C���P�x)�.�3zsfqk���OD��<�'�O�%�b����?)�����


�A���ůLLi� ��$[>���(Ov�?��ia��<��O�u��>����� 96�R��Tp�ٙ�o�i*Q� F%.����r��<1Yw��5���;�>���T�Ifo>g>jS".�(�Q@4�T��?�`�1�Ya���?Y��?Q����&J|(-ά(�*���GJ �R������O����Op��攟��'xL7M�t�J	�fD��A�|�p�Sv�qmک 5DI"��h�~��r�j��
�cT/�Z5_O���O?���V�$=Dq �(�'���4�����1E��r�'���'\��FL!^[�Ӄ6>$q� <(���b���Y�ȗ������O.�$���c>�.�$�O�]�NK( Tb��O��*�m��=bN�o�MR��r?iG+יqJ�sGt�4bϣ5���E�%,���N�ar�5p��A��?a����B�������F��'�����]DJQ��O���fd��/G�i�bm-GH��2w��OF���O&�Ĩ<!Gk	KK���?���W�^@3�џH��ҳE��%3�� `���'%�I��M��ix��1�'��`����=
�	Di��g04d �m��
�	̓C�6�b�	���x܀�K�x��dͧ�?��S�y)�4م�!e����F ij��e��O��D�O��`"�)o�X����D�Or� {��8�RAY�~�tJ�I/a�z��p�re;���O��d�O8��J�UE�I�<��IÆJ�bDC��˔�Hd�!�&F-^����_$�M�c�:ň�dӽ]I΀ϓ+�F$ӱcq�ݸT��k茼�5��\v|B��_�!1#�^������Q3�M:�?����?	�'i(H�H�	;�^��EŪ�:H�w�
�����R%B�qS��O��D�O&�iX�|��O� �0�ܣ=���A
�y�)�c�<�P�i �7"}C�d�';9h�R�O��􈜓n�D�H�<Clp���@�J��<�g�
/��`�'�UPH�� �b\������T(�)������40@�ւ~���������	�����$�'�>�i4�����E�G����&@���E�*����'eR�T��$�<)%�i�7��
]ނ��CA�Е����AX�M7e�0���N�*8��Dӛi�(�\wM��F��<�\wo�]f� !"��R�\�@�KR�e�.y��M(���$�OT����t�q$�I�O�4�E��V���f/۷P���<A�L�K��,��I����矘*�ǻ�,pǀ�)�`�7앁�J��-��d���y+(fӬ���Mڠ$C<϶�+P�'��k�ƞ H� jçן����Q�2P� O�O"i��Wy��O`a"��0ZF�d�OR��OIp"Ƨ@*�4C�V'Y���$�O�ʓx�xx;� �?����?��'
���
4D2L�He:�&xi��G����'?���M�4�H?���C�L���2Kn�#��-�E+CA& ���r��=�L��`�U���I��C����T񡌀���T�-*�����	2�IN�[I<]�I�T�ؕ�
��x�������ğ�'�̵Z�Fd��H!�?�������/0�Q���'��'�"���d�<�e�iY`Ģ%
�|�L��ALТqݠ(�6of�T툐*\1V�󵃃�L�󤕚���R[w�Ny�&��pJ5��9L���)�c��7z�q�)Zߦ��a��2u�ў�?����?��'N�@�ɟ� `(��`V�<�i� LQ�Ab�]p#Ï7�h��S�����?�2 K4����y��End�V�^D��+҄�48���iլ��'�Vt��TD�Te�����O�}���g�P���E�Y3�'&Np��� ��h!#$�[~��Oܜ��hH5H���Ǿ`Pı&��	�<�b��G�E^�d�ON���OH�?Z5��J�����O�0��d�5��3���+pH$8��	�OX�sW�� �'��7J���p�����KЋ;4�t��3o�=\�Z�����Z�?O�YP���5��u���Ɔ{C����	?ž�ӡ��s
�8��Z����G�<�?���?I�GXT���L~���?a�'m�iQeG܀8|-���^1f;f�{�r8jm�3�����O��$ÒwS���<�7#�K�z\�",ٿ'�8@;�	L_qxu�&���M��d�HU|�رo��0�͓|R�If�s��X�5RiP��$��@�o�2=J9hwi�ty��O�Y��]�O���D�Ol���N��S�<6�Py�D�&��2+�P�6��<�Gm �c*O��d�����4�~�D�s-6����v�~ܡ,Ɛ{`v˓����n�d�@�O@�j7����iV�{pU�K�/#�d!DfKbx��.�(@� 3O~��@����y¥�4���?�B�/.�� @@ �^�5� G\<zpJ�[$@2�?���?I��?I)O��0!�bV�:�����~�x��P�|H�F�'���'+x��O�˓U>�փg�L��W���1��Iy5+�$�Д���	:�H���*,�X1.�Oxu�Ê��u��ʉ-����u'�r�ł%(��1��p���a_n��d
��a��O�D�O���MV����N�!�� �l�QĴl'̝&-�����O~�dC5@��}�Bi�<I���?�%O�{?��s���h�)�� � �W7_;���\)��p �O����U��Mid�IX@�d�>�\��cNR� �2����dq6��F9�?Y�"_���?��bV�ሥB��?	��X1�=���^'�գ��9D��0��?�)O�I��L7c���?q��zX~�SC�4�Ҵ��xx��s��	���<��?��WQ?���#"���-D%Ҧ�[2b@�t	�
H�DS��D�g�!s�b=E��a݅����O�ɓ�QXy�A��,�I�e��m���^�S����D�B� ��O���O*�d�O�˓#\j�ˇb�;�2�1�A�Z�x�@�/^�p(.����?���?	�lq~���8�I?�B���Å*e���H0D��oڈb(b�㡉�,6.���k����	��F�g��3�O��b�l Qr�EIg��D�X؀ش!�r��r�#��'<��'���+ݘ}��w���9��P5h亱�� �n�1ԉ�G�D�O2�d��Q���<y��y7nH�bJ �)rH�2�ε�`R�y�ViӎZ��O�2an�4��iP�3qd���� �I���ǧK�(a�Tn �~�����Ort�d��?���*':副�?���P�ޤ�0��
�vD#�/��h�t[R�,>9X���?����?�*O"تb!�24��O ��
�3�6�c�)��.J��!g�x�&�DÙ)�Ijy��l�R�l��N��7Jz�q&�ȚT`ؼ҂�Y�(hm�LR�a[>��E)y�a�F���6�Z�k�6OP��!|��DL0�E���6r��J5�	--*�zdnJ��?y��?��O�o.8�HK~����?!�'��9��tB���Վ]V̌����H��H;���O@����T���<�$�	Z�����%
���D���9� UK���Ms���&nBP�1I��ZV��dgh�q�I��2�D�aG�-��Q`���:�\!\����._��1p��8�?1��?��' ����Ǎ�#t@���ʿ`z�့k
���Dڝ�2�8���O��D�O:�)�BP�˓.5� �N�;t|���l_H�:*O��lZ��M�楞c?�S��,r��\n�EY �K>J"d��Ra��R�NH���G8%� �4G��<	u�]+g�l���n���'R������E�0j�(p6pp�"mX��R����J
P���O
���O$��<vm-� ���_�cUÎ-^��C��ʣPi�Ov�d�O.e*�����'�67���E�4MB(!�R�k$E�=C��2��27I@H�T/N41�b�#m�<S�� ��n)^L�#+��]�;d�D��.IV�t=Bԯ�,;�x:�BX�f��x�����	�?���I�Sԟ�K��9""�è1l�<d'CTy�'�,��W�]�Ub�'�2�'�4�'KX�1W	�T��5���B�J9Ҁ��Df?�!g�+Il���4�B�`�B����� ���?�a��|�ʤS�˃�(@�q�FI�)<����?� C�=��I��?y��״�~�����?���*p�����bF,��D��9�D����?�(Ohl`�ݞt2����O<�$A!�����TCAlO2`� �8����s�F˓���I���S�49�� ��9b�PV��?����L�^1c��T�.�R��@
�R�|;�,��6��*�e�쭻M���	�%��l�,O����;P���w��N���Ƶ��50,����?9���?����?Q.OH�@j[�=�n�v�
�TTJ���/��%w�U�dg�O����O�����z&�	ky��}��ՃCf	B��Ș�m��er�q��� ���I@�@�`�֑BT;e�8��I�r���q������7�y���y��9%�˒kV��P�o�)>~�� �O�Zu��4Z���Or����pVI=�⢞��,�B���`��Q��G���tx2��x�I������dT�̖'�6���Æ��J���I�7K.%���O�6MS�t��$��h=H40�O���"�2E',%{R��zl� F̄0<��n����'d^s�!��<��*,��$�Ɵ`)6��|vvD���~�4=�'`�9R��[B�J�y���������󟰕'�rU!�c��X���'�Ү�$r8Xa�F�[8h�fD�:�"�ڣ���+?����M[��f?!e*ڝ$%�I	��8��[e�Ý�n`��d]ӟ�.w��0[�b?0�y�6OFם7�^牶h,�@kb�ҕY�<��.D�)B�U*R�'�?!���?�n�2���@M~���?�'��B��g8���L�*�d4����!� N�$�?���?��� ��}�'
��:=Z��q��\.vLqt!�?�l���;g�\7���^`������?t��� �=OPh{�4�u_c�䅋m���&l�!,Q3LD@4��g��G� ��F
7�	�	��P�	�?W�b�? � ��ǰ]���9T�ۀ��D#d]��r��Lﮝ�I������?Q0nz>]�ɪyu
 ��ʘ�x��ȩ�U�y�� �'�7M�m�'&�����+¬������0a�I3>��S�ۿ.\blB�!#�|�C�����p�.z�I�^��_�d���`�que^2Z�ބ1��ĄhHUr����M��B���?����?����䏉y¶!cP+�O.͉��7(�(x���!+�N�0 !�O����O������p�'��7�ͦ��D��|3v��n�ى�B;��y�ac�:y�|��" Tן�8@n]!��n�"@����'+뮂�;�D0L@*��b�L0?V��D�U�iSef�ן���ӟ��S��, %?Y�	0=��i4��+&0N��C�9b�Z��Iޟ��I�M����E�ݟ��I��I�+d��0m%,�`�eJ.@����$�����!�O���b�\�6-�,���.@[�	�:O�p�F��hB�*lܧ� �X���D ��u%\�YA\��"�7kD�{�B�'�?I��?�4�L�"�hZ�O6H���2�L�%�?�����$�!Sv�=T��O(���OT�i�0\nԨҪ��>�2�ήIN���࣠<),OF�oZ��M��!�Q?q�b>���Sy"bpr�ǀ	 �)�7Dòt�7B�"`Q`�śd���k�uk�(�O$4+�zy""&h5bQ`�a �0`2���1���DTvDPx"��O��d�O��d�O|����$j
vN0#ĉ�ne� H�..��x��?���?YPo
\~�R�,�ߴW�^)�G�>D�h���/���� �i�� ��t�D G���y���@^��;9��� ��?ͪ4a�r�ƹ9��ƢF���d��������� �ޟl��՟t�������O����̐�	n �	��7�iE�IFU2����?�����o�q�T�'���� ��D����qy���@Z�6�Uܦ���)������<v���P�L%�r�J9�CDY'� (��aݘ.�F�z����lz&˝�I��ؼa��ʓ����9�4�r��'�>e[6�Q$�zD��FV�Q��٠��'2��'L"_����h�( �	�����mKn	�r�Ѹq�&� ᄗ}nڴ��J7����d���4����	��l�u�>���1�Lן8;�i�r�F�ϓ4��"��W�qU�����F�T��?���1(�T�Irď{DVQY0	H�d�M���.��*���p�'���(S+PK�Z��/	!]�ʑi�����H����?����?���@�'���	+/!86��98��򓪚!%�;��YH��6B�o�a� �V� ݳ�;O,��vAQ��u�d��qod����� N<�d�Gf���(L�耔'&��dL/(2Œ"�4�2��e���ݚ�L�z}��@0��rAXʓ����Đ5�?q���?)��Z���O�ډ���a�z���K#!i��su�����榩y�`ˉ�?��F�i4�'O�`�۠n��@d��Pjݖ=�':�ƽh����<�� �J��02#
��'�v��+x��%)V Ӽ=)T�V�a�>���D )az�V��"}�7�'�Ĝ���ʠ#!�\`��/8�4*$�'���'�u��O�˓����j���9T��%k
����<3[$��f:� ��#�
=�(��2O���ɥ�u���/}E�\�O�L��	x�N�� N؍!Y���ǎ>V ����ĵn(1O����STQ��PҎt���"NO��\�A��O,���Otlh2Εt�˧�?��sİ�=�
��G؁v��(��J�[�����I;�?��iE�/�ĩ�ݴ�R�b2���`I��<Y��A�y��9��M��f"���>�����/�O^���NIy��Oh�P#N2^1O�j��՛6��P��X�Ц�Z��1�	q�ʥ�篔�����P��
'����$��b�eA�@�W/0�F_y2T��ش��f�X�C��$H�����O<�|��L�*����� �6�D�) �Էv�Dl[�j̑q�L�Γ�u�޽�?1�J���ɷy��"�j�I��y"��2R���K�c����!O��?9���?����?!-OP�� �\��H�
�m@��Q�ܕN��r �O����O��.r���ay��w�2�1Se�],��0g!
l��x+�-�ߦm8�f�T�(��4&\H+J�	�Sr�A#���&��e	K*����O*T�R��Tg����c�=�M���'�A��L>FV��'��O�<�� �?q#�ЃNDdĲ�$7?��x�6i��J��a��#�<A���慙�|���?�w?���l��gd�!��ƿ)),��ųi�7�5?����w�И�̟��3�m
KU�sv�(6��`{��ҝ>��Dk� �4.6��䎑k�͉�*��(PwY�p@�qinQ	҆���?�b�07	�ɹ�M�?!`�I���;�?I���?�������U>X��d�OZ���O��!��Ⱦ}f]2	�t0~�v*�OVU������'+(6́��)��a��lBp�H��<)b+,1�N��5Hg,t�ɀ;O�pQÎ��6	&��.�哄^��Y01WtL�C*�,D[(H�G�y��Ap�A
�?y��?�&�3!&!JK~���?y�'{���cZ�|�,�Q�/�AX�f���l���?����?���6y�'��d�:'����a2N"�5���S7��Af��.��7�9[
@Pi� �u���ZF1OL��&�u��b���S�KN%��E9 �"R�r$��hOy�j�O楋���3���OT���pS�G�'`��Y��`V. �Iq�oЃ]��z��Y��X+�?����?��'V��Χ�?�g-яZ�Az��J<V��A#̎?��d�O7MM���$Ǧc~�ap̟T���Ȥ9*R(�"I�2��6��v�4H�3DöH����i}d�?�s�J�� �?Av�S+^^���F��@���k"B2P.*�?A���?I��?�.O\py�B����d��$>��.�qF���F�M�jl��$�Oh��L��dy¡aӞ�o��TהMZ�S�^�Æ�$s��\)C�Gٖ!Xℕ0u�L�I�D�"zW��i��������d�����B��!�t����������ٟ��ǟ��xr8�%?��I<9�@�K]=u��\�C��0AITE�������5�Rܛd�dy��'�2�K*�~2�H`>ܥ�Rǚ�S<�C-N�6`�)��}s�aS	�M{��1F�@�ڠ^���I�UL��ˠ풆t&I8�ř-x��X��Z����;�\ʓJҤ��O^��� �'.��'4� &4`�'Z��8�� �!Dh�)b�'8�\�l�s�9\���I����?��� �#fXA�L)��m�r���	��'f�7�����C`���Q�#ʦ.�i�,m��ɰ�h8�a�,��W>��6���3����L��yR��J$���'tz$j��<��(ڰj����%�O�<D�q��;_r��3�W�'���')��'��I�Ox�0�U�K��`��MO�!"�2U�iz��I����I���/z�h�Ij~2�'���{�����` �4���0l1�i=���R��<-*G�_x��ܺ�嬻O��m�``{����ٶ]�����&��dڄ����K	�-�T�׏�?����?�'o�Bd�͟�����R���p�1ȝ�A��4��B����H�'���'n�$lH�����'��6��QC+ʂm� ��m���P����O�6�'��䌏.8�2T�O=�4͔2�R���c�h��;�
5kXqQ�j �ml<,`�'�l(F��<QS��!��D�ܟ[�	;����ɡ/��0;�$W:���u�Ѣ	������(�	蟐�'��pׁ��T�r�'y�H��iGR��e�9� ,s�/��R�ݡ�y"�'��I��M� �i�"p��'冰j2B�[�b[T䕷,����	U�i���G��xS�kךH�P5+A�XF��ί�y���)-n}����|+4��8z���D��O����O�B�n|�䒟l���O��	�c�z�B��$+
6 x�M#O+��$�? 
��/Vr�'I��'�`��'l"4OֹQB�ԊJ] ��HGXh�tm��H֐��'`��y��&G�:�ss��gu�q���X�5���8g���σ$E������@y�	��O��I�}���fL��������� 1��{��߻Q���78:�F�	Iy,(8.��W�''b�'����Ӿ����'䜱1 ��2�����L�"�*� ����������@Š��"�(O J�����t, 4�4d�*�i#�AS���@��,{��y�T��MB30q� #�~ʓv��&-}����h߇��e�6�riV���)�����I֟t�	sy"�B1��x��'�8p��n
q�<Q�s� [:�\���'���'u�t�'bb^��{�4]u��âQ�)��,[�Zζ�C�%��>K���� G�Nс0�Y��y҄Y�Mq��;S{���%�|*35�:��`�U4�<p�F4���.�I ����'��'z���־ �OO��z������2Z���C���A�2�'DRa�ƣ����D�O:�dŤ��d�{�"�{b�V9ui�kBg�{]f�B�'h|(�v*�$�?��'i�ޱYr�܁v�6�Γ-SV�N��[�,�v��R����'���(�~�dϺl��1�'�������u����?I���?�fز$��Q�biA$z"<�ۦD>�?����y��� �?q��?��'V�Z����+J[���Q�H2FATi��׀��d�<i���?��e�m?yE�ՈKQ��#/�:ȳ_���c%ô�)��C=�L�wER�=1y�<O4�ݔ���$ήC/�9�'�8lxF��P�z���
�*������O�H!�)N�o�@�d�O���Oz��<iR���P�!K�.�{G#��.��Q�2�ñ��$�O����*���xy�'�I�4`N�={n�3�왽P��'�'�4Qe߰�ç�U�yR�\olѯ�A���Q��?10��ʉ�θ��C�!̘Y�{�B�	1�x�T��b�rp�j
�R�C�ɵ&��akދ}j�lqC���'k*{��м���x��!x����%Ŀ	$v��iۅaRȌ�¦��3Cz�; ����ԣO[4.	��%%[6aja!��G!�b��xͨ�����*��U�JG^�+��/1sf���c3FT��`RkK�F3J�ȣH�UL`��d[,��4�!�&�Ti�F9R|�5��hL�Z:1�"M�}�CaP�qYת7����mV�~�X���n� ��
ۓ �* �ȺR���avƔ.z�N�h��|�܋�n
pKYm��_��i��ͰN��p��œ n�hZ�j�� $��u 5I߄�A���L�{g�ÄRz 3��ʌ8dXk�B˼i@���"?U��|���X6��;��~B��bG�%ٰ��%�
(	��ͻQO��M3���?	��`d�h�^��PW�`����^�&�e?uD���x��Ç�ܟ&���OV^���Iɟ�K���E�¸��[-p�*����⟄�ɿf����Oe�=O���K��4wD�`|�9��Ji��2uV���0��j��ݟ<�	�d�'��LҀ�̠oP����y((!�l��WP��%�6���?���O?�ޟ<�	��� (�!��Dܠ$���R���&��4�I֟��'��+B��@�Qǡ̓܆D  �mŘ��7�'T�#�'�b�N��~���?�������1�ҥ�NO�-љ��Ώ ��9�/O~���O��Ŀ<�%.F�M
����`���z��ƟXV�X�L����	�!P��"�����O�ѻ��������GE�gc�P�C6f�2�' "V��jI�����O~�D�)r���/!�
Is��3%�r��"��`?y'�C؟,���d�n��?њw{#	#�����>72�)w��?�(O���j�����ş��	�?�;�O$ ���-K�,]Ʌ�R
�L�R������O.�{7%$�F���O+V����AQ2u�V�L�]�̱�杻"�i���'�2�O����$]�Q��HT)�z�����I?|�D��(�����H����O��1�1Y��O�mt�AЋ���>6-�O����O���G}�&���y�'୰��J�1j�1�6΄+`�X�[� L�0��O������O����O�Hq��M7�\��1'P������O��$\AȒH�'�d)Ҝ'`�F1�~�w'�{���w���rEX�"���-O�ua�h+���O����O�ʓcS\�	a����Н�RG\5�F���X�t��ɕ��	�(kV���i�O"��1Q�`��GpId���(Q=�P ��&/�$�O���Oz�l��t6�O<E�b��?��U�ia����?�rn��<�&�
���?��I��L:'��<�5C���5q��}�fl�E�Ey��'��'�I�qT���O|	� �p;R�ͧm^��fڒ}%���!�'5���~�iB���4�����O�韕��$�����veka@[�F�2�'��[��P�	����'�?ɝw�h�*uC�(3+�U�Z2�F��F�V?Y&��hyR�O�����9OJu
V�	:�6��ㅂBf�HC�O�ʓ`��(��i��SƟ����� \�X� S�хX��N�@= �3�Z�4��
��@�)�S��������Oʈ"�"�.�q�B���n7�6m�O����O���Ty�o��|�@'K�"Zb��#�tE�(��`��?1�# �?���S��O,<xR�
d��`�+��u0u��O����O����io�˓FQ`�ͧ�y���<E���`�Ho��8�I�:#lX8��'��$�$~�h�D��dk�� ��LZ �C��O���X5���f����'�yrF�Y?�;l��PvHɫd��@��(2��&�|�`<?9��?i����$ٿE-v�ED�:�!Y!��,E8lZ`yb���?��hP�,�O��ɴLW`x���[�yM��w앟g�f��	̟��'��'R������rWF�
�XM����HXt�W�Y�<і��ğ���ID�&?�O��bغҼ�X0.˅w�J #��/$��'��P�L�	K�ėO�b؛@�����	1D���D��esB=O-8�' ������)>m`�!3��s��Y_�$��*���x�����?a)O+�iz@A_>�����H̻?�r,rċ�"5V�&�L���p�I2��O��������"*�.0�FͻV����m��H�Isy�E�K��7��|.�M��'.��Ɋ�0ɨ%����X(6k̫Y�!�$�<��T��?��S����	S>,�d(7�Q�x�:���gʀ!��D���n���O����OJ�ɶ<�r�T�|"���7�v���j�R�Хˑd�;�yң��gRHMEx��4�'p�A�F���{8���ET�:��B�}Ә��O��H��X��'88���'&�#��"�<�xA�U�DH]�d�mL�HG�'��'%��HF����':��'�dt��!�^p꣯\<'	Aّ�'�b�L�� ���̓�?��D�<�wl*��pJ��a�&X�䬜����?)���<���?9��?����򤎯�����(��3Ĕ!��L�]9<Y�2�j}��y��'&����'��4�'��DRBd*�� #5������[��j�Od�$�OP�d�O�ʓQg����O��<����<EVؙg��+c��<������?��-�<����?���;����@�8�IR�٤3P�6h���N`�	ܟ��	ݟ�Ify2BT�V����y��Xn���c�O�&�^��%�F�?����`I͓]��e���?��I�<����yB�4}舳�G� �ۄ'��?I��?*O(�`�_���'�r�O&��#]�)�n�K�"��m�Zɺ�k��y�IВP,b�'�JxJ�O\ʓ�yg��S6�����[ܦ���]�?1-O�j���������I�?-˯OL�㑫B�v�Ji��j��;�jq�i�lY(���O��t5O"�Ģ<A@��K�i ��LApă$�~(�5�	�d�r��,t�:6��O����O��	�G}2��y"H�������e���l�5�rl�5�y��'��	-0lb>��	;_j�8b�_�R�2(c���-�ߴ�?����?!Ǜ�y��Iy���IៀK@L�M���ū`��B��I�3�D�	埸�'[�������'��'������"b�����[:�@��'JZF$8 D_���GAt���%k �	ڼ�5	H!n>��*��u.^4��[yr��y��'n��'���'��	��V���F�96��jq��.Q	V�H�Ρ����%<���O(�X�1Oz�I�O��$^�`eFw����ڑx��Lc�8O���?y��?�+O�p*�n�?zf��)� ���ЂO�aȲ�O�5�7O��R/e5����"���O���9O��� U�	>F�↎�1[N��7$�OT�D�O��D�O��vD)�TT?A��*,���aC̔�V�@ ��m)s��������P2x��RpΟ���T�Z���̓D$l����Yʒ\�F	ˍ
�	�Iş8��Ey�l�+�D�'�?�Ǧm�S�z��s$�/��	H'$L�!P�u�k����(�����Ib�P�3��uޱ:���~���aa�-l��Y@��O˓Q�N�t�i�R�'���Ox��G��1a#�.�r�k��T���Θ��?���8��Ex�ꃜ�����E&/'���#"B� ���d�o���n�D��П��S��DӼC��DJ�	����	��p�vժ��?B|l�O�&�(���(�	ß��Ш�F�p�s#�Q�n� ��(���M���?a�f�Ԅq�Q���Ih���I�h\��ǁ<_���S�Ufx�X#���m�@Td��<���?���y�
Y5A��ZU ��(G�#Nm����?������.$v��	ԟ�8�j���;G�l���.&mZy(��c>t��'�|�0�'�؟��	՟\�'�0�Z�n������  Z�����LW�k@�PQ�p��?���<�'�?I�e��)�V�t\�5��LMv|VA�j��<Q���?���?a����ć>LiT�I�'b ��:�Ht33l��1��"!�y��'�ֱ��'.���'�c�*�y�BO>~G��@���P�m��m�b�'8��'��\�P�C���	x�i�#!�����dҶ�дb�OH�ʧ{��D�s_����O�p��9O��4�����E	�gj�i�k�*C�^%�c,�O0�d�OT���Qu\?����,���-\f<�AG� T2����GAD م�}��i7����7a�����di�i�6�B%���H6�׺̬#�"�O.ʓ5�����i&��'�R�O'�듋� �\�gF@��H�øU0�T�Aa�'g��'y�̂�'�'�=8J?i��G_1��\Y�nZ�L��9ւ�O^��&&զ��I�T���?帪O�1B >O�ɉ"'�;%���It�\� ��O �QQ6O���<���\̧�?A�i�=8,�1O	�/���ǋ
����'4��'Ȩ�C�<��˟��I�Vl4�C�j���A����a�*��`�Y��%�`b��Vr��ş,����ܹ23-Ղ���^: ު�c
�(���d�D*O:�a���U�4 ����O�X��w	 :J!��E mI�d��V���a��D�<����?A����ň{�z�N�F�n$R�L��| �c��`y"#��<	�H ��O+�'�h�y4�$X�V�V����AjPb̦aRr_�x�Iǟ�%?��DX3�����<�\�A eʊh�B�(1��<�DEi�(���e�hY�Os��'s6��s�'w:�i�&\� �ҁkS�Ģ��s�V�4��ğ��I[yb� �@�N�ޜ¢ň�I�4��LǑd�Js`�ON��B8]'�dL�lrb�',̽��{�VD�z��5&�L@��'��?���?i*O��}��՟$��(��Q �MۊnGf�X��Ðz�ʩ�Q,���zA��O��dU�F��%�de����`8Im��J_I�����Oʓ?d��p�i3�������򄘈9��PUj��"T�#�O�5 ���A�'��#T��y2�|ˍ ��S�	I꘨ੀ"wR>�sAJԽ��$�5{!�%n蟌��@�� ��*gB4H�x�ɓ���ecSJ_�lb/Z��|�� ��Oi«ckt�ܑ�u�*�0�f�3[<6�O��d�O��AmTGy��F�<y�Y�r B�Υwh�}p��Y�J�Dը���?IO>ٰ�����?!��?q��� ��0�ț�w�	��Ì�?��;"��GW�8�׮�O��ĝ� ���<*���D�����֍J"y�y�' ����|"�'4��'L�Ɋj#�Wz#��SV,�%0Ap1O��(�>˓>�F��0+wb4����?qs�اc1��
c�]�q�j �A���IX$)3������O���O��0���س�OǲĲvCݸu�r�h��oľ ��'�i��?yƪ�,��I�O���'	���D�7N�1��JF�f!b�+�#SF��?q���?-OԀ9�'K}��!O��˴ȋ#3`��*qjӂYD���	�|䈷����@�O
��ǩ!&f��!?�ϖU"
��)�v�C�aR���������'A0��#-5�I�O4�IE?WE��(�`P/Jyd�	pI�&�tP��O�l�5�'Srn�8C�|�4��բQ�E�thB���<PŰ��'�I��:�Zݴ��)�O��)	jy��V�]'�x��H��!�Q��a ����?)�C�4�?�O>����|�IJ~�u ��	�Q���*`C'.2mV>P9b�'3�'_���'�r�ʔ���CI�on�]b�f�*~0\�E[
+�������Q���I�O�L����gd���Aw� ��������0�ɕ5:�\�.O� ��O7B쒏���ś7e`���޾-b�4�d�Nw�CE�<���?���o�9S"�@�@7$C������?��ɝ��=m���O�-ئ�O����v4����\5�P
�mƢT�'����O��$�O��D�O����.���p��a�d����A�X�˧D�O���V�=f`���O�4���O��'L󄝍c��(2u���`�S�@?��fW���D�O��d�OLʓ�&s��OhPU/�	`�SL�X�L���'�ҵ���?�G��� �$�?�d��B�z����|U[T"�<����?���?)�%��	8,���䌺��8򡃗ea�����2	����OX�S��ON؃`�'��O/�� O�H����)t�\� �5e�J푠��O,���OZ˓&BNa�v��d�'���B���$A�r�Z��:F�����CBg?�u��̟4�I�:�#<�w� ������"4$�`�!=P�P`r����d���XoZR�d�'L�D��<I P�Ml��Cdj
m*�E��L��A�	�����g.�tx4�O�t�#H��>���2掰w��� u�'Zb9��kӈ��O(�D��nt�'�@���a���T�ʬ7������>=�-Q�@�4Ex2��;��'*�+�
-�L�sJS3)8�
J�x�$6��OL�D�O�`2�IDyRe�8�?��,���+� �;�(���:9@R�Ì��' ,��y��'Eb7O��D���
�2��i��*m �'^Zp�@0X��2�o>���$
���韪����͠>L�Y�/P[��Y���(�ď�$w�I؟��	ԟ��'����	ްwi�xbPƎ��nH̈��/O v�'0r�Я����Ob�I�� ���@JXt�zBc�0�4���ן���ny�e�O����^��Z�{�CA%P��՚F)�t9��]�v=�'�2��S>��I��j����['�ǣd�F=;��%t�:�de�<���?a���dǗ��]&>�� @��d��N�=p�4�V��ӟD���%}x���"���O�<#����Ǫ�P
/�ع�D��T�m:iN�c���:s��9BC��9��3f`�?G�ݓ�H���j�;l��XqNe0�'Q�h:�����?a)O���0��O2�d�O�OB$�dM@�a�fm��߃�f� gM�O�y�@�O����OB�O����	.�)ƽI�i"�K�<^�N��wɕ9�V�'E���O��'�)�7��$�O����^����E�V�*_�d���8��v��{D�'�(ق��N�k���2��R2@����'����T(��(�b�Q�L���[�k�K��(���}���� ˿+����Ɍ98�$@y��X 3�,i	�׀ >aL��t�ؐm_�[d�Ѡi�X��\�#�I�;�.���� �J� -�ĤhT�OL���!k�D�x����܈P<�m"�]6H�x�A�&%�V�U��$e��!tp!�	џ �I����]^�������v�:�
�78�n8s�� m	�I4/�j}�u!�x��g�ND���#B@�	�(P��]��e-���";�8t㇉_A���'��:���B!��"l'!A!Rk)?������_���Ӵ�ՙ&OlEh��q#1�Lh<����4�T��V$�6J|�R��~��%.����t��'#n
Ua^n����,�P�`tC0&ӢD���T�'���'s�j�	w��};G�'��)�~8d� �x/������r����5/�	����$������$!dL0H6��ez��dlE�w	����ހt\D��[y����$ D|���`�-�;� ����bX��*���O �=��<u��<��`Y�,s2hХ���Z��yҍ6�I&+�(9�M�)*�(S��X�~���'��)8�'��I�5C4��b�n����ئ�ʃ��kh�$�m_�+t��B�V��?�MX�fbh���?ɃF��a{�x�k!E��ӺC��8L��1�m��yz &�j�'��C+��Z���y��?��͞	�n%�3싵s=�ܻS(j�'�J���?yH|r�ɢfQ����-Ym���¬d��6�O( {�Oҫ(�������ꦵr�|r�8�S�$%·�?Q���1��H��@��q�q �.5'剜OLB	ZC$����	t��˒�X
2�iQ���eɠ�Lɘ$��L-����O�@�c��j��s���l��3$P��L�H�%�іR���#�'JԒ�6��>�W+�	����
�)�rAs��&=���2 �ӽ\ΚUh㌘"*V��i��<�I��ڴ�?��	!������"oW�8� �Z�7���?���hO�Ө=��"���Tx��Y>�⟰ҝ'�TL9��y�T�O�$��8J�<c�B��D�0�R��(��2�OF�2�M�M���aD�w��"O�÷kØH��1��ӣz��Q!��{�(���˝$��d	$>����R�ذm^)ʄ�2n!�DvƝ�""XJ�Ѣ�f�?T�!���[ ,�*_e�N��%�$G�!�$�U\��S��PL��,Þ�<�!�ˑy3��(�j��f�b� a�	�!�D�*h�|��!9}��<:f���!��<g|	��a���ܺS.�6�!�$�\�8\	��	�z�LH��M
��!���`z�<�D�[��\�p�C1,�!�$��2�bh �F�{��QpK�!�$�Ta<4�u,^�;p����J�	�!����r�͑gF]����"GT!��׷.o2�B��)��j�!2!�$�.V���$F9{�5l�:�!�$X�A�1C��^i��u�l8lY���9M�����2T��J��B)�y�e� �����К'�re�T�yr�D�(�T誅L�;<���cI��y����I����!F��r�s���y�"<g&4:�D�z#��#;�\]K�'�Z�"�Y�N�,)��ZC�<	`�I�k�2$	�/� g�z�&�YQ�<�R �,��}
��Ȣyu�i�Q��R�<a3�L�N���6�T��l�a��H�<e��5un��"'��+&��8�CK�<a�F��2ʾ�{2� k��] '�F�<1��Γ"��b��L�h\�P*�~�<9*�[5�IQ���N�m�v�t�<�`˼e��Ɗڃ�!�
�y�<ɢ��h��ps���0z وO{�<�n-���!�G�7! ��h2&/T�4{ ¨�yB�C���$�7;D��ˑ�C<L6�-Xr�Q�2�a��;D�� g�3P��y�#���L�b -D��(�F� Ϯ0[� _#c�[FK7D�б6���:j�%��E�
!D��JD��|xr`�Z�8���� <D�� ���4˘�8�� R�V�lm�u�#"O(�3�EY��0�cBY<D��r�"O܍��Mчw=+ը5CY���C"O��(�KQ�cZ�Y�fڐ9|2xz�"O�i�l��v�Hq ��dk0mI'"OrU� �ʃUW�2�� �2X,%A�"O���3��?f�V$�̠lE`�2"O<cC#�@�`Y{�%��`G�م"O(ɰ���ZE��-�.Y��l��"O��I��[):�m�v-�&m��X��"OF�:�ev�S��4�*y����`�!�$Y8Y����_�m��9%E��Q�az��Q6oh���2Z�̙`�'z��-!��+6+�!��l }���ȇx�>2��L�)��'�:�".+��(D�d���B�Aa��0�0�!�*Ә�y98���Cfj@�*��b�'V�H�c��yB���[�,c?ObU��ƕ^XT]���튰��O*l;�o(8��qE��W8�HԫΘ0�2�҃�P�S0����Z�lPFb�0�&i֣��G@ay�,om<}R솲#��d�*H�i(@�[2I�T,qE/G!�d�1>��q����t���uK�a3�8���J�悐��2b�zX���F-Ƙ��@�n~FB��'�zyz5D-*���9��I6 >L���V&UA��N�}K�9����'I�)��2Od*�ˑ")�.,1�LS�a'\�c�Ot�E"I,��N�l:�Q`Z�)*@�Ib�Ә��!��1������'C8�=i�A�6�R X� �<5,&����±&��5h�I�L�%����J�x���d�ّ��H�Ұ���}���1f=�O�H�#��#c��l�&�U4zl�d��\�f�(o8��jDiڝiy��*��l�ʔ����l��n\�}��d)'bI� ��������y�g�!iZ�PW�O�J��e���V�ZtB���i�$��[�5����k/�i[92�銔;��͡Ao�7��|�� RB
-ɆO�ݑ��
x���p㪃�.v�0�̿&�Ĕ�'��4�>6�N�%	����dR�����UN_�P�O�]�0
��|#��4��(�6�Y�a����L&"�X�������@�Y�^^�\C��??�\1��UOP�U���I�e���ۃj�-%V��U�|"��S�X(���j�S/@,��t�.�'�Z�ppH_���YΓtX���dȎ=�i���F��Q�,H3���U�,(��H#TnY��O�8p�̕/R(PUC&)�sru�����sp
}��X>�PuM�u=�vhKCp�+�-PL|L�h�B|�3AO�j����G�Q���cUh&k�"�y�.ңٞX%9�$ݤE�)#�j2�Š��ֆ4��mB�`;���B�ɓ�#1=���5B���y�#T�'��@��F4�h)��� I;H�p�`�
�pt#PM�Lk���T�$6��ɳfu&��@R�\��"���-�C�ɳ8��Qb*L�M�tX:��[ZB���%����	�$ �-���ԔyA����4xl�B�_�m��R�w��x�%�{��M0���={X���EĞf��x�/�W��ⴢϹ4��58� �4������E^Hi��>��� �cF�%yly�.F!1>���b�*J	z��V���
}T�j�k7Qf��%�A��0��O<H�ɴaÚRj�(��P�k@$���#��L2���� �Y���Cy�'L�$tc�O���ϗI�쬚��Ύ8����W
O@22"��CiF� �&ܘ���OD*��i��:�M����>���h%��[���GI+���!h4(�֡��I!%�d�lơ��I�A�}:�oX*:.���6+�6@ѰB䉌h�| ��$�V�Ȑi�� ����P��� > `�OR�1�#���h����O��r�(7����>j��<�р�JڸD�R�i�m^xw�h�&O�1��㞰{��OX�g���9����� HK|��G�����U�]�p�b ��V�e���+�EC0�X���I'�!�� �ED�8��n�(��0�`U���#�%Se�Bs��s�D��+�C`*��'5n�^�"O��P ���o�.�R֦��N�0��CP�t+a��0��h��'[�h#a��c�0�%�%GR^��J���X��
�h�]�'	�ZP��M(
l����;4��s�"D�B3�y{D'X	&���sQ"ғ#�*Ѣ�#Ѹ���F�� �ON�a��KO�I�Mz���if�t:��� p�j��ݸ#�l\�7��bЭ"U�i/\�[�d�o�n�o�u�BA���J��5�,֓h$�тFB�Tbn� B� �y��>}�P`C�!�"\a<��1�=<���G�7$5�eC,�j�����)шbd¶�VçH��W�}���B*��>��$�C.d㰣Z0<Q0[S M=AiŰ�M��
 ca���g(|O0M`� !b�\���D��q��I�X0�'����TH�>kzh��8��ؚ�����ִ*3e�);?�B�I�Q�i�S"[3c���FX�|0xb��9�l��^X���S��(� ��B7r�0֫��^B�I�A>���ק�4_8Rd�@�W�WSX�H$�y��:}%%�g}B��+}T��
Ì ��9�e�$�yrһX\xD�׉����#L��MkWK�M�.1*�:|O��r�L�T:= �@Ȋ��e#��'�i���o�-�	#�4�uD�r���Vւi:C�ɔ���R�IC<Â��Uh�W�㟨��A
6+7R�E��\�&�F��ׇ)���5�$�yˍ�6���AA�ͫ���ZE�
��ذyc-M\�S��y� S��Zh���j�2�����yr�_�L��jB#gtZt�ޒLV�q��{rO	f���$�.ڬ+�皗A��U��&�%`�a{"ռ+� �'/r����M�5��ɒ�2���o��	�XaqPX��ٲ!/U�]k��E�M�z��m/�&X9�����֟����F(2}����nz�i��|�6�8!�׽V��0�B7Fk!��@'2��[B
Q&a��Q�`�9hS��?%�m
��\jn��C��3���d���3��Uٳ.N�:E(HgJ-Ah (�"Ol��POזkr�9J5�ۚ?^��7fF��jUɖ��US��٣Eнdh���V�/9�	�)�JL�FJ�1'�X4R��6-��zRl	!�LȺ��4~���%��|��ᚶ�T�p�1C�	vVL��,j�B�1 '>lO(	I�i�o�X�v�ʷW��z��6]��Amґ%��M�FkU,e-�T�%O-�.�;A\�I�$]Bjʵ���	S����z�>�1��-�
���$P�����7lR�0�8�j�n 8KE��1*�9~�2�)3�#�4�0�y��ܕi8}�@�#o?�g��y2�\!p�\����/�h�����6��!���}.�L�R(�[��LK� t�H��B�TܓgT�%z��n���(ql�/2���I7[�t� �&��,��/��)��l��̕�F�-�H��c	,��T�E�M��L�1`�'�8,�@ �	 �t�����J��s�{�V$j����A� lB(P�$��rS|y�HފMQȢ �^����͌2�j�c[E�<11���*/���M(L@��$�΁����.R�Ф���Q�'Deb�Jܹ(,ޒ�\I�;i�L�P���9��ԭ�P�R��/D�0�K $(�@� J>J�-��-0y�0%� "������ kך��p�e��|����J8�4��D$�O���@��l�xu盱/l>�pR�S�<�  ���H�T|�=��&S�&�>��d
\�F'ȸ.#x@� Ы;џx �#먤���F�C�x� #�����9��A�wQ�h��"O�<CΖt�r�
�n-�:]8�P�`�1�H�B+�̪��?������ }m�c1&S���e��C�6x��C�	�@��#�Ы}"�PBEI'���1D�? u��I�$P��A�O8�3�&:��d�pET�_������C���C��&;���	��ޱH���QH�*xC>�H�BX"]�	�T�L��p���<ra�����<5@���7XR��d���� U�>�(dA�'7���KQ	bn�-R%�{�~�r�']�a�bǋ� D�!L�}$�a2O>	G�|'�m"��=�R.��Ҁ
:Mr�X�N�U,��ȓc��8�j�$l��`8ClA�<j��3��YJܓ5~̣|�'Ulz2�Gm��8��߯`AV�S�'v!vi t2�,�t���Q{�'����6)�0n�Bs)\|�P���'8�Q����:_�bܰB	޲v���B�'*����i>�|1­j2����'�V9���Q#g���A�;���'��������o{���FY�2tY��'^�d��S��lx@4��*�
�'�00ѡ��O����aץ?�|Z�' Pt�f+@�j��Hc�R6c������ b-��J���PXy��E�pn��B�"OXQ��뛔*�$���W�#ڸۄ"Oz��f�0����l͚1��`"O��صc
Z���p�I<�|y�"O(	 �M�#�=�@�+�,e�`"O������5��p&�_���2�"O��BO̓YW$�	FӬ? q�s"O ��Q�;U��Z�gʦk�9�"OX��+L�O�ʽX'ѨB$r8:r"O����j�ɢ�����|2r��"OvP���בa9��#��)y"(Z7"O�{�✈qo�Ũ7d �G��0�"O�5�v�Y�@���2����t"O|$;VB_�!�:����U�f�(�"O�lq ��7�`L؂�>?��)ʂ"O� SVgK@L9r��"Ph�!�"Oz���i�+� ��̈S96�"O�����ڸqF&���W9`J�"O6M
���?)Jpa�Pm��6����"O�U#�&�F�*�=h��"O�$���²e���a��K-sO~E
�"OT��W����ۃ'U4B(N��"O�@���7���0��F6z����"Or�r��(���M�.'�n4�"O\�,D�a�Py���)�8��"Oz���$F{����Q�!�pԘP"O�mڗ.��c^��h��5
��"O��a��H�.:-e)�#;��<z"O�B�����&�ޝ�����"O��+aŎ�Q��b�j�u����"O'�:�$ B��9�B�!ll�;���"TF<<Z��<|OXi"Rf��B��1�Vh[�*�^���"O�01Q�
3��"v�P3"���a�"O|���hN1,�\�K�$ڭ.+��K�"Of-���Ff��EW=`(� ��"O�A�����4y&i�r�ɕ~'�h��"O&a��M�2�0�p�J��� �"OBT(`�E3/P���Rc�I�h�@$"O �"L�0���95b�2m:9ۗ"O�Pk�%M�n���k���?;�X���"O��X����`��Ϳ��U`�"O��T�%>վ�C��
r"O�=��НQ�&�Ҧ��0�ڀ��"On�x��|��uX�`P�W�.]��"O�(0@	6i��q��� R
Ԁ�"O�@��ñDtd	��	PX��"O���GF�%uW�qC��B��cU"O�J��E":�hdI��խ�;�"O�ɚ���-~?�ܘ���d�<���"O�8�4�A;���JC�J���"O�l3��X��p�ڡh/A �"O6�^:��'-��B�����c�)Y�!��?k����E�)Nc�r���!�!��L�Tcv5+qD�|^��eEc�!���A�����-�����!�X"*�1#1��k���Ӓ�X�!�dŸNM\su���T}�!{uY}�!�DC�%��EhՆ��g��`��X�:�!��@%ll��	?[b@j!NK�+�!�$�;X���R�γ(<m�-��A{!�$�<J�E�H��Y�q�SL�Q~!�Zi/�=# �U��(�*(Xy!��)v�����v���S�U!�dA�E֨��N�Pd0z�)C�!�� �EC���r�j�OJ&��%�"O�y�A�>!��3 Ό�:�J�0�
O���p��~�q@4B�j���`tÙM�P�g�@+����%yd,؃�HR6Y(8$g�O�'��� M�t�� ��;��[�&���Y3G���[����p���ȓbA�k��P(��;��Q�S�H(�O@�����D�`��l`�OAf�"�
E�^(�O?բ�P�'��1�+Y�p�D$�:7c��2���J1@��'�ƙYcE�S�g�	U�l6�.��!�M���0Q%`<����#'Q�V��6rҀ�!��j!�G�H�7.��)�',�O��K�T,��y� �D
I2|� �'M���f��!4�傩���0d��7�jU3Dǭ*]z (��6D�L��L�$s�X�mĩ:N���5}2@ڊW}��Wo���p�~�rA�#sQH}��˅Q�N��.Df�<�a%®�B��ҿ��Ls� �^2�Zl�>�g��9 �>�O�1�҉XmKp�x�����%�PxB�K%n�vp����5_��9CG��4]�졆m%-�zy�->�Of�  �Q<4�*��0��.��|C!�'����p��.^Ī��s��4�	>\�"��X6!v��ye�%D��x�+���:�6�׹K�y0��"}Rm�w1�4��L�'h�~b'�G�C��*dƖ�6��D@fd��<y�ќE�Ĭ`K{Q���)Ħc� �$L�>�b��L)&�>�O`x��
��0�^��j9���^_(<��L������^��U���_�d%�@`L#%T��u�'�6YQ#H��L���K�)D\���}�
�w��I�@\� E�X?�'��a�-q�p�#�N�-[J������L0*�Ы���,9�P!�����'g�"}�'�d`���B$j"d���aJ*�ڼ��'�A����+^���A%� ]q��4lZ����*�OTH �S^%~H�ǂ��K2L���'�Hq�I�ky���R��5�p"�([�N8�m^'�y�Z�!�� ����Sp հ��A���'x���@���?�s��i �j�kX�o��,x�d&D�����8�,5�v��.4�.m[������$�L�'�g~��� W�D�,��Q�0�$�Ϩ�y �=�j 1 .��sԒ�J��K�`H�����}"�*�:T;��]�c����
��0=S.���@a-O�C�A�0NN�Qp��M�}�̘S�"O���A'�f	�"�j���h��$�n���(EM0�'T�\ Z�#�L�81R'+K�%#,�ȓ^�������ER�A��)�@U�5����PuF��O�*#H[4��B��;�x��"O��0�E�:���aF.Pv����jًkL9�"�OQ��M  �ޑ����,��<�V"O�-��+X:siv�s�O�c����s"Op���+Zx�͡"�� [N��"O,�#��@���� \8&�u�0ȃ8ukPnQjX��:��V�-@��F)K���+��.LOb$�%ʏF�5�'��QàK�P����]. Undp�'��E�� ,3ҝ��咽~g$��y哿zo4,�e-<�<O��CB��>���3n���Ld��n<r�h2힣"ϊ$@���n*�`�F#��"���'�D�����6mG�*��Y"h�@��p7�*D��s�Y�L����/*Q���[ѯI8#"�e�TOН)��|r	lI>X"-�m*�$Gϔ�0=���4�x!�#g��l����1d��]K�OF�b_Ԅ�q�1D��aVE� s�0�7X�]��I�F2�b]Q?]��
(ZI�� ��r
���!1D�4�5K_��$� L�� ��c'�$D����G_5rs�)@3$@�ߌ�a��"D�<�v��,0z���-���Z�1w�!?Y��Zx��Q�/�%�Ԣ4�ׁ,�N�Z@2�Ot����O�*�����c�� ���.�9v!��z� �S�^ D�}8�G@+Sq��@�π^�π B��wMH{��9��-s��0F"O�y� 'J�� @�UT����3O��4o)�)�'NJ����Iμ�c��*{�(�ȓ~��1$�1&����S�Ċ��x�'D��KG�'�e���ļ-Sv�s&��Z��d��b�AZ��k&�9��(ҟB�NВ�-L*lU�؇�e5ꍹ��P1l�J(
�!Y)e�P�G}ңߚ�h��������I�e%�U�D�(�O�5�cb�>��q�PF8�R�ٴ�B�	))���!�t�T�Ƿp������:3�⟀ipɃ/&:�Ls�fÕ(���2�'D��f.�.T��eɂ�_�$@�{�+&?������L�����K����n�11r"OjɁt
��=A$�yM�#�x�!�D�!���D3sy���`�֜�x��.hV!�D	1wq������ԓ@��'�$b��04�h�S�I-�Z�)��߻]&hIק'D���.\6O��R��9���,*D�@C0�J8�xHp4fҁR���GI5D�D�$ß�o�n�Sp�N7>�:`��6D�L)��ηP�5I�OK? :L��3D���]�2b~#�a]�Z �q ��0D�<)�'��kFk_
Ǯ�/D��ȥj��	t�ժ��� 4P!�$-D��2�����p����>�ؓ�/D����-����DtG�*��2q�*D���!Q�g ��φ>�|@�'D�H��&%�f!��ʒ�
z.��u�9D����DC0O[,-�r�0
>��pD2D������0X�!_ ���/D��bT\5g�jA�"K»7R�� gA-D��2�Ń/����%��L�̬�&�5D�|�Q&����z�I��\f�%2\O�TRb*6�$��Z�:�k�^5����ɱ1u!�$�=� -:3d��J��X�%8qO3�G$�)���+,��s����t}�\ٱ�ȧ`!��/1-�f̖6mP��s&]/�~���(�$E0K>��E�ŭQh��F�/T\���Ɠ(~� Q�!ưr ��0T̉RV����"��(�5�O��K� ���{�GF�i� �a�'����*��	9kl�8�oc4H�f�tQ�B�	�GchX��\�:��I�۔nej�OZ�J�ä���x��i�=�\{���3\�Nġ�+�h!�$S:{Q�����:d_�Q#Ƅ
iҲ����\�D�9u$�?�'�^����Q(O��ѐ��KPa]*�'q>9:3B��EK��F�j��Š#J��S㤨B�%I�t��|2*�#s���B�(S��(pJ7Ø�0<I!k'Y"��C�K�yd�̓T�py�B�W�<�D-L�!N��ʓy꬀�ۜ(>��U��5:�Y��� 󧔅��uy�,Wm�O]�RNӒ>�&�B��K�n��0b�'G8u��I{��yQ6K�5xryv�K7?_�᳙'s�Y��+ϡ��Ϙ'-�hȇ,�?kю�����TV��'�r�j޺Y~��0㌏�`}���\1if��S�)k��|��)f���!7A�)��R@����<�Eb�J��"���~��,�6�2��H)m��#��˜�y�Cxj��ʚŸ���$ؘ'8���8/�?����D'`���h��H���k�B5D��0��V�`�� ف��K�i:s��O��D��O>mi�O%�ȼZ� W�Hr�E��"O����![Et�!�M�,_]8�s�"O�����{|�i wL�)Wx�i�"Oڔ�Gm(���j�6s���"OdmPG�_zGH��`i]�@�ZQ�"OƑR�9b�|��΋�A��ٲ6"O� �I�Rk�K�`!�E���̈C"O�z��ӠE<<���˘0�4��"O%����jHQ�˫rt�p��"Or``�Ɖ^�Qxg	�i��E"OVx���	H��
�'׿9��0�"OD���΂�O�8ǅ)ٰ�q�"O\��-��{6D�efǗp�Z�5"Ot��5�P��8����F���H�"On(:���38�L1*���s~^�ڕ"Ox1"�9S��hR�V�Y�2<�"O�0�-_\M������1Z�����"O�]�&�G�!R����u@�"O����&Z�D�� bҁ_�\� =��"O�HL ]��ȑ�C�b��p�"OJtQՄ-���B�>Kvv *�"Ot��Ԁ�:s���b�(4l�l�"Oz����^ľu:�KX�A9Nq�"OYj��z-d}�uT	 ��H�"O���<.�
稁�z���C"Op0�2ET�~�:�E�D:Ӑ"O ��E�#T��u�$��'B���"Ohw��(s6V�b��N\|p1"Oh��GD0Fڤ$�(ۿ?�9��"O��QS�DZIŨ@
V�1A"OTyWc� d��J�%u�
Ԛ"O8��ȅ-"KU��j*!�"O���X�E>�(z�j@76����"O��AQ�I�}\X �iS��H�"O�����@�;A�$hFg>_c�]��"OxP����u�c&�t��3�"O43G��6�R�xH ��"OR5�O��xc�ly�#Z>Pz���"O0h
Ղ��KB��aA?	ΙI"Oh�Rg�C�^ݼd��A�4[����"O�4p�� s�-��O>j�H���"O�ɢƊC�pi��C䪔�e��$"O�qx�M��,i��Z W���U"O�-`1B�47�ah��T6$ ��"O��#N�-�jt����6�V��b"O�(y�CO�f���ier�G"O�%a����<�����{bX)�"O�Ԛl�aW�� q��3m��[�"O���ɬH$���dE�yQ����"O�ĉ��M?hz�I�$K�^9��"ONM�6j��6�)r�ɿ?��X�"O��k��V͚�����Д��"O؍r��� LP�u�!�xZ��"O�4�v�M�5���V�ͧ'K��y"M^6V��(�v��=^��Qpm��y�n59�䉘g��#Hl�,��ݑ�y��D�\�s�&݉+`h�i7���yRH��#�p�a���%���u�Z4�y"�D�J�Z�)��V6 ֶ}S��/�yb-D�i�rLx�'�yx�-j���yrJ�
Z)�]���j����e�^��y2�V�������.v�a1%�Q��yr�__�͐�S#y�� :�.ۑ�yB@
�{$ƁY�@�<^T$��cܗ�y2���:S�͂�C74E�\���Q�yRc�-r��̀";�z!ó�ۅ�yRA�VRPr��>B:���^��t�ȓc䠡"kW�G.Xӆ�UZY��~d@̚��՟<<���^�8ɇ�U�:I)թ�1h�Nؠ��	cs$��S�? &!�^�wF�{��5(A�y��"O*1��M�n[J����ɲMZ�9� "O�|ҰÉ+��	��O�W, 1S"O4%Xω/B�8j�ߺ7"yW"O�T���_�_��kè�K��)p"O�)hRF�*/	��g�Y��+4"O2��.Y#�T���hſ>�,\�e"O���2GZ�j��Z�╍[nN�5"Oz�ѩ��IF�����[T����"O�B�X�o&5���J6�\P"OΕp��^/��a�1�ۯcf��D"O���H;+�~=�Cg�o�Q*3"O��+ .�x���#C�t2�"O��rL������4�*?����"O<0�m��^g��� 	�Bz���"O���gʒI����V8Tv���"O���-Z�8����uh�q""O|msW%mP���?WxTyZ�"O>A�A	��d�)���c��"O��6��#���*ÌK�'4��""O�H����*�N\�0��v1��ɧ"O��8Zݴh�V�:e�t"O�yʰ�r jL`�F_]�pX3�"O^\)sg�#���pL�1%�P)1�"O֝ �a�Q�B%���g�tԪ2"O�e���'(zi���r�jP��"O\	�̜5.�T��B��H�t0��"Oֽ��	,4,�ĳ"�9���"O��3p���J �_�L�U�j�<I4 أsV�+Fg����w���<��"�*kO�� �a�X-"��|�<ɠ�Ջ~��ᖂ��3�.Z#��{�<��iԕ(�V	���ڼ	��p�a�<9b�ۯ]��(f-��vH�L�FNWH�<A�K�+ER�`���V]K6"�]�<i��-�*MS��_@@�%g[q�<i�KY�n�H��({����Me�<A��8+-���e'X5��qM|�<A�v3�i��J$�^9Z@k�|�<a���-�A��kO� x(pl�{�<	'�X��d��{ϲ�
�u�<ᄧ��w�n�Z��M8�z��׉�n�<Q��Y&E��s,T�h�5c�Ei�<�0��&Ɩ�pH�7-���8�IN�<	ɛ-NL4�a�8�@�(�DN�<�`��Q`\Y �պ���WaF~�<9�ME5���Qamķ%&��`*Ky�<��EL���`H��)��`"�A��<�֡_8����f"5� T���p�<��b^�ɖ�A��9,�>��AE�l�<QA��0k� ECA<,���D�	R�<���ss�\�n7By^�Kq��t�<���ĵs��g+-B�����OY�<� �,w��Y5D�)a�T�5�^I�<A�B�7:�� $(@78i���@�<9W�U(f�d���	M�Ν��HV�<�q���ȉY�E�,�p��U�<7��$�`P	6�C��d�b��Zw�<I%N�	'�z����M�er�<ys���HH�`Ԛn�����@x�<ɀB��jj.��2��)0�yr��t�<a�])W�&� �l�'uj����
t�<)�M�	H���C�C
T|�R�T�<�A)�7x������Z�Yur	C�	RQ�<� d��+o)Fq�u�vΘ-20"O�d8�+h�� ǩ�
-V��"O��Y� ���o�]xU"OZ� u��wa��7��_��6"O ��mP�v�݈V]�t�Q"Oj1�Wa�IE���0�N<P��&"OZ��S�ٱ-~�8��J�����"O��I����}�I�k���tȒ"Oru�b�-�=3Ƥ��7�z�8�"O<4��;K�$Mi�E�=�l��"Oz�K�,�S�n����*4"O�]ʲ��N-t=�4&���!u"Oԩ;��5վ���d]�����"O&�!��O�0ܔ�cP�A�����"O�D�u��u�-�塕�J��t�"O�Š����3A8,A@��7_�
	� "O���@/«{�X0{ F��v�(b"O���'��O��Uҗ��|����"O T��l5VnB��_��C����y�Cǰ#D:��j��z�1�b	�y"�>SjV%��gG�a���G��y�+����!R�����`�����y"
�cA��	��FtW�J�(T/�y��U�x=j���ǅ�����D�y��/,�P��+�5�h���i��y�&�)<0�0�I�J4l��V(ߕ�yb(ʻme洰�`DA!�]��K%�y�g�C��1�ڸ3���B׬�y"�؅�����eY($�2أ�#�4�yIW�_I`( �W!H�Y@���y�h��Xq���I1H��hV���y¢W8�"�S�#�U��A�)��y�ɞ#)�LѢ�*?^鹷��y�K��$d��;������y�ហ�X�����*-��w�Z��yB�Q0D�=��b��ʑ�����y"�
"���4�Ϟ_fHq����yb&���R�0]*��ȕ�y2l�5B�)��$E��z����y��7Y��1��2T����ї�y��@Dh� +B�.Eؒ!���y�J��'W8[ �l:>m R��.�y� �G�����Є-������0�y�O�-��2���?;�	D`�0>�I>�DN�7#?l\*F����.8�7T�\p��D�i���f�1HN�0��>D��{�H����<�B�}�p��
(D��b� Ao����0!�W��(Z�2D��х�Ʌ&��\�S%�%`j���.D��`�cL&2ˮEӦ)ڱ�H��2D��yg��~�x�D�Y�/���Zr�4D��ږ�L�'>�\��J�'V�|��C.5D��� �Y���E��<(F���'D���テ*7d�1v�ܕLX��2D���bĜ"��p!��2< ��w�,D�ı��=[��I���̺7��0{g(,D�� T�Y8)�������.��@J��&D�T��f�3,��`��F�W�ز!$D�Sї2P�����M�Ʈ7D��BP�F�W����@AҀ9�Gj(D��B`�׋g�<A7'�W0 1�'D��c�!�	��@&���}K��8D�P0�
ͼ� �s�.Qđҕ�+D�LY$�2��[�N0Wn����*D�� zy���q{�n�=�~���"O�� �%�3^�*�kG�H�@a"O�5�o�0LQ��;�̳Ab���"Of�Z��ByQ���3�x�S"OH��a��q���(ҧgLH���"O���e��=J��01aN	W�H�"O:$r� ��"�B�Y����,6N�zc"Ov��#�f�����&P>t5R���"O<q
�(��+���SCG/N'h�7"O:���3�T��!�v1h�kQ"O�d�[j���癕F�\Z6⑍�y¬͚t�|!D&	0��@v�<�yb�y��!�ƪ�� �h��%���yb�L�PS��C�%G�X���A�,�y�oܓ	&�M���?86��4�Q�yHۃC��	�%��7����ӅV��yR(�4A��c�Щ/GT}3t-Ǯ�yR��^���`��+, ()�ì�y�%O�$�%B�	-!Y��7��yrC׾^��2ꀅa|�1��7�y�����a�,֩S�
�#����y�ɑ�ldp�ˑ
Sj�Y� �y�AU�`HZ�@`X�OA��(@ 	�yr���d��PB�K7`��r ���ybk�"T��0�S�_4kA�1B'���y�*Vf��J��1o��ᅉ��y�吓 �vlx�]�1�"<�p��1�yri@9`�kl�-�d������y�E߭U?�H!����w
$ � ֗�y2Ó�B�w�J�rδ!�R��
�y"+����F��*h,E�'��)�y��R�X�Y��ս]��& G<�y�ʏ�IEQ����`9���d��y�K(n�X�*V�,Wx�U۠m��y2���Rtrt�UA��鈠��9�yR�	�(�Հ\�
J�x ��ܗ�yR�˄SW��r!��o���Y ��2�yҁ��G%�, 5�Çdd� �.N��y��	ˬ��4���B�A�R�B�I2@Mp��i��Ve	�Il{�C�� F��Cf-��IeH-;Mɮw~�C�I{G�Y�ԭ��,^>%32��9!�nB�ɍ[ �ġ,Z�ۤb�*|%8B�	�h1R!���%��HX�,�%�*B�ɨǒ (u�Ӭ=��Q�)NкB�	�.�ĸq��fi`��FI����C�I7u��@����[�^�����W�C�ɯ7b� ���H-2>�5QDG
��C�!y���R�<J14�ssBR�B�Ʉq(�K!�]�f3��e���2��B䉕Y� �!���_�h;�� ��B�I�K���u�F�@���7ӾXLlC���-��LG/ ۤqt�ҺN�@C䉱C���"
�cc��@����@�C�I��d���8'
bq��F��2��B�16���ٞ:����CM���B�ɪz�|	bJ! Ȩ�!�bG�VC�Gf�-#�A<m��U#�%�=�B䉗���
�`^�-{�
w_"B�ɬv��y1�DV�"Π�����k�C��n]b'�!f��I���W"�B䉝���x��°{Q�9�`��/�C�	0J��=9a�1\�� ����[ZC�I�d�a�fު�xM��bW�.�XC�)� ����E�;UН"v��U�8�p"Ob�j��H�N�k��\�JV��8"OԠ��^����eŵsQ�#�"O��ЀX�p+��|��y��"O`�Rb�F�I�	�%	��b� �@1"Oظ��(���� �W�P�la�"O�\kS�(S7>2���B���"O.���&�R�wmy�`}��"O��!�o�?eU�P�򅘸w���"Ob2'�ğ-X�`���F2U����"OX*�6T4�A�D�qX `96"ON�Gh YM�d�,�� "OZ�#��G*2f�!����nr����"O�@0l�(5��eʣ�Ϥj�Zkf"OH��'\�	r��:q'Z P��uj!"O���C�[�����6E^�D"O\̸p�75�|c�c0~&�[�"O��pg�U�Q�����$i��#"Od���c5_ƅ0ea��%��08�"O���E+L����@C"��k� ]`�"Oqq��j8ny
q#�����!"O��Eʞ7�,�r�/�R��"Oj)�½��K���c��
�"O����#�4A$$���~��T�d"O�Q#ӆR,M��,3�i��	t�ؓ��O��=E��A��ƴ	�I��Pq�ĝ�!���d�.�¢�|�|H��#��!򤖯NIX�D(8���yL��6�!��x`�zO�,�4���I��^�!���<s܄�(e���H9����HF-2�!��(O��pʕ��7����V��!�d�i�1{��Ak������<(p	�'�D��dF#
z*����	v	Dq�O�=E�LC/��H��c��)���O��y⁔1 ��$�+T���f���yR G�}}��Y��q�(xHӋ�4�y����7�x8�mPY�|\r,��yrჂ5d�"K�N'�,��B���y��P�7�,�kƯZZ�,��ğ��y���z�ؽ{�!Vd̄��IK/�y���{��k�Ӝl70`�C(�/�y�M�?Y�,`ŢE�Z&d)cFC�
�y"j�,%>���D4@3�h0�yb'�D�v����hЃF>�yB	N�Tz���!�6{������y��L=�R0+r$I�m{�y�F�J>�y2D߂J,(A1ɆY���R�-�y��Q?lJ��'�L]B��ө�'�yRC�+*�����#P/MTҰ0$,Ô�yfC3�T�ׁ�:G"<�뤅W��y2c#��	�oAA���ISd	�yB�G�c��m@��PS�u�2k���yR#ZrJ���&ޅD� �A�l���y��N��E葤Ll���0bAW��y�T�4qZ�"���"p1��A�9�y���`�����5	�/��y�瘟Nla��M�#	��
A˃<�y򄌁Cô���k��V�T��p@޾�y"o<|�h�f�"G��`E]8�y�ξ8�YfgՅp4I�P+Ţ�yr�-O����Go�(q�(T��L�y§��B����'p�be�&� �y2�U_v�<��d>_�����#�y�_\�l�a�D���L�tG�y
� ����<�q�s-OM>�Z�"O��k䠝�ud����Cے[G"OV0��B��[��p�)���|[e"O�a�RM)) \�i�k��$@�i(ў"~nڇ��- �LU�4���*ә��C�I,B��Aؓ0�Y�Оs_�B�I4[�v��e��	���.�b1�C�5DF�A;v]�G��T�q��%Q�C�IP0�eCO�.7�8��,Q�y(C�8s��Q�rJߕu��`:��{��C䉉c�6����³�	{1m�+��B�I�d�f��	�/�˂�ж���'pa}�`��R00Y���~���lВ�y�A�UK2�jf�~t��q�"�yZ���PfŁ���(�`I�n��ȓ��,���U�K�Ri���F��ȓm����J��6��q��o�{�x�ȓ��I�d��>b�L�����W�V��j���F	�5!�	���l�E�ȓ�y��Ŕ}��,�F��:$@�ȓHؼ�h��IDL	����/�ȱ�ȓM����i��RoT�bg��p�l}�ȓ+�4[��|��	�O@9丆ȓL�� ȖX�|.��iq�Ǽ`zPl��~�.���F��f�(��ƈ/�i�ȓC�RYG�_)Lh� x5��0W2Ʉ�N_b9��#^�Pi��"K*~�>���쭰��H�!p��iڨ�`�ȓ8�Y���>ఀ{')�!a���Ji,��g�8fb�8���7;�ɇȓ<łM�Ee��K5�����#y�����Y�1��ŴeM^��A��  �P�ȓt��"�,ҠU6���B�n����W��Q�WE�Oz�)�W�P[M�M�ȓz�ɪ��T����`ɍP��E��ȍ�d)�I@N�
>�v���(5k6������M�;f�`��l'���3j�}e"r�� _��I�L����C,\������Kpm����=�^�d�⵪ͷL�L��ȓ4�dy����p���^z̄ȓ%�n�{0�W u�"D!h�~�u��Sl^pC��]4Ih���"g�(�������%X}QtѲ�CI�Vq�ȓ^O aˤ�.3�\�yS$[C��,�ȓ.��8P��ėGU�p�� �Z���bu�pR(D_>-�vE�p� T���t�"��7��" M�"d�ƅ��S���7�1D�nHZ樌#�%�+D��{��22o�d����r�q�	6D��.ޠ	���¡��м��4D�`�1�$}��k�C72��
�(D�P ddF)m|l
@,`BJ�Hq(D�4�"�]�}TĖ���@�H�5+!��GChT�舙 )�g�F!�D�@_F���$i��]�e���!�$ܟZP�D�����k�0S)CQ !�L�pY�H1&��N�v�"v(�!"E!�8Ҍ�%�[��n�´f�FA!�� O|`;��n��P#b��h�!���*�Q��ʔ 蘸[���]�!�d��)�Qy��^�N�"�:6��� "O�� &	�`V5�I��+���k�"O����$C<@$
+�nݼ>�uhw"O� �q�5�4��عp���9w��"O �ò_��@H鰨�f�.��3"O�Q�&d	z��@�Οn��8@�"O*�HG��`f�,I�AM��Q�GL~�<���'Q%v�`V�
˾�*���O�<9&�M3*]�B���\��'	H�<�Sj��l�^5��IZ�V-�*�@F�<A�D¦/���3=O:��S�M�<� �}I��@�E?�I�N̊k�pC�'q��%X��@�O��y�	�(�C�Im(2��V�П��q
 I
dSpC�I�k���ӳ�M O~5�V"�6 �C��X�Z�#e6
"\M��Pg�C�	P��u���XqY���*�=?��B�I.�N���e@T�..FJ�B�ɶ<Z`�H����}�F%��K��B��X���J¨8����l���nC�	�,����7������OjPC�	�,�)�Fְ٤P974$��B�**E�,��GʌFIvH1��^x��B䉍|5�$ϧl�d�pwaG%=�B�	�%@RX��,'T��H ȃ�W��C䉛ld�Յ�$g���r�Ł9Wg�C�I�ePE����6@�:ĀF��]��C�	�Q����Yn�e�l��!+�C�8y(��ٞ���UK��tB�I{+l)�CiӪ-���lO�r�nB�ɑEF޹r ,T-N��G�M�dB�	����x��U8I`� �A^2HB䉍,u�R��F�Ġ��&MB�I�"RRH��%�k]�A��.G��C�I �����I!��)�%�7�B�I5,^���猋:�(!bf	hnB�I$#�V���%$3@�fH��>w~B�KS� k�W�Y�1��!r�JB�ɗ(~���>^hʁzC#�!q�0B�	"�Ђ�S�0�L��(�<6p�C�	�yw�-��D�ee�T�H���C䉱n�& ҢPv�8�oQ<aapB�>4�
l��#�''lܬU��7o�,C�rC��c�!��f��BŌ��C�I�3�`�*'b@#DB>0)6��k�B����[�b��,K �����+=x�B�ɴ[<�2�,~���"ʋWZ�B䉋L^NH�6�C��B�PBD<yK�B�I�6b�-2�,D�4��Cm��C�I�@�q�GQ�G�"���ƨQ�C�I�PV2i8�jŶ[�
�k�aŏR�RC�� 61�d�r���=��A��8'�fB�	I"Ab�H\�4����e���C�I)t��%��b׮8fV�*(D_8C�Ih6�<	p ʿ{���R�����C�I%g�:�I�(
~����%K�{��C�I�}#��"�c�\�j�`!�Q>b�!�ߊ$�8��"�� 6\kBdǑW!�č�%��L���ɩO�.m��ߎD�!��(�+F%P�k�<U�s�K7!�ă:��D�ע@(���4�	�]�!��v"@�0N�6�8AB�A�sv!�D��}7��ǨA}�> KP/Ɍj!򤗮^�x�g�>U�u@"@�@;!�9H�"cAU�g���y�IOg!�Pb�~����ךe���iͩT	!�D��1����Q�(��L�W�p!�� bZBEU�����&�*b�95"Od]�$)ځqݺhs�%�~�N|�"O��Э�!Q�0��$A�G��9"O�<�u,K�5\��J�*�|����"O�a�5̨����� ���"O�*��K�ةz�("_:9`�"O�͊`W�}��� ����"O�)��ǋ^��Y1g݄�V��"O��0".T���Č��Q�`%�""O�������GY�XN��u` D��#DO;R%���3�Xl	��;D�LX`e_:4(��2i���d!o=D��;u��<ℸ�@D9T��1�?D�@P�Oݗ ����ŊU�F���7D��1�g�IF`9�壀�e��t�5D�\� ˓��Q�� .f�qР@3D����dZ)w�P!�k$�5��6D��J@	�6B�t�oP��!�*2D�C�ȒI�9�K�C�L\{P*=D�`��J5�"@�G�_}1V �46D�����%�A��$���L8D��x�$�$`dvI`�� z����2D����aX
f��H�#r|"��7/3D��X���S;�SMH��m��/D��I�&�(>RSC���A��@�-D�l����3!P,����>	�r��G?D��j��/sCz��g'ըI��Hń>D�x�Gg�'�V�h6��3��l{7�&D���Y�BO>@ O�� I�/:D�8��	�p}��"	�%ju�����9D��)W�%�F ��%B�r a<D�ISHS)"�ZW�=�r9Y�)7D��KR�� \�
��Ǳ'BJ±�:D��a���7��bwa�4������7D�XA�fH�GI�@$^7�h���6D�̒���Is�$���ޏTSz���2D��c6-�rӈ�ˇ��m�R��§4D�d�"�A�ZU��)�OV�)z8l���$D�� ��E(.��T���J��dK#D���ď�OΜ�Ƥ^ K��t��<D�ܨ����	G�ǋa�`�Bj'D��2���t�������q�|#E/ D����Q96�4�Y��]�y[��PP�!D�x�`�q�]n��z�p� D�L��N^�CJ�L�v�t�9
@�=D��*��Ke��E36LK�d	�e��.D�( q�ؽRa`�)�ʎ0�N�+ŭ,D�HT��P�2��4N�Yd|YX��8D�0���,�ָP��ܵ�l���h)D����Hj�!�
�#out:��<D�܉���,_�К�U	Alv��(>D��`'�	���Y�o��;������'D����bV�+ц���C��aG2�r�G9D�\��(�}2ģb�0�pĒ�,#D��c��7���p�.۱� �p�� D������	8��[1`F?iԨ(6�"D�\��*B�
��P�&��`��K-D��8 �N>6�����iu���E1D�h!��g6f�itF$���J#�-D�X���� C6�1	#p �tZaf/D��[#��d0� �v
D�@�#��(D����O���XC��æ`���z��%D��R)�>�:�Q��@�ИTh� 0D�ēìgH8��ىMPHPp�!D�� ���֒�Nxza)V�Ojn�)�"O�d�S�_.T9!��G,!yb��W"O���i\f�@q�°fv�Z�"O(��q��2f�P@�b -dL=��"O�����Ps�-r�lZG.RT��"O�)q�F�%J"�Qfܞ3�$1�"O����̛� 4,�4�B$9&�=�&"Olm��՞F�>hR���Р�6!�䙷g�p ���S�>�V쪖��'ay!�dT�E�I(�K?$�BDx�l��!��f �|�ǎH�4S��sᬑ�!�d�
Z�n��u�ˠ_��� ��R�1�!�$؅50�����xT���闺Q�!�5k�0v� ^\Z��h�*�!�X{yȀ:��ڿ>�T�����@�!����L���/
��^��dFɺm!�H����ڂ��1q똄�&�]A!�9g����� '<LY�4��8�!�ĉ4i��0����2R3 �#�K�B�!�d��>��<�B�E2�����G�!��-F�Ijy��I3@�.y!��ץ� 5*u`�\�x�UΖD�!�����O�9�p�ԬO��!��;?��"CU��H��ʙ)0�!�D��z�bI��!ܱ������*g�!�X2�J4�(X0m�h�6�Z�-�!��/˰=Cu�E�����B@Ú�!��Ҁ�R���7�L��n� K�!�U!ߺL���l�健hA�$o!�dԓa��a:b� f�y�J �!�$�B(z|�䤓�`��l�CL��w�!��ۗP���%5��}��kW�P�!�d�6���KհU�K�e_�h�!�D�]���rBH�N�:��҆�d�!���s�x
0��'�T@��F� �!�d۟� P*���n�H[a�X�>�!�ěX4��Gm�#Xy�s�_1!�E�a�f�)Dƃ'��X
� ��>�!�D̳xR0�eT�m������d}!�d��8�^D $��Rr58�ܳv�!��:2�B�BD��!*U�w
�-�!�H�^M*���f"���b��3�!�$D�Vb��Q�W ���m�.n!�dP!h�\h�BI�B���+����!�D�&ljEccÆp<ޅ8S�\�f�!�$�(8��0�I��F*~�8*ն�!�V5���	qAɶ"%Ұ���Ry��@���� � s��xG��Dp� �ȓ\���	DZ/̢��eN��q��	kyr�'�v�ڇL˷a�|�[�@Q�y�����'���J_�����
�Y(J{��]��yr�$P�Q2P�Q�P`rd�rDЪ�y" ӵ$-��6.��Y7��!�yS�D9Q� 0/�6}�f욲�yB�@�_�\$�@��#�$9!�'�/�y"���e��4�PC�O�<�xaO�+�x��'c�Q��#�v���8vd�"���۟��?����(h�� |oԛ�^�<G�� ���A���̃�j�x�<9��k$�q#�d�>lP�-H0ˁK�<�'�v�D�"wC�Vdx��<�ҠA� �n 0��6PN Lx��o�<���ϖlߺ��e���{ZpX� �p�<�6 �0IZ��ɵJ��UCg`�.�?I���'�2�'�ɧ� �@�v��a~�[�I?pƾm�s"Oz��5,H8TBHy&F� G��*�"O8��0��6�R=Y�$�5++�ͪ!"OR��
�1	pp:3$��f���S�"O�i@�k��9fA	����"O4٠@�D4r�c��<	O�D�A<b���X���ݠ����H��l�'�j8��I)��dX��UNSB���'#��k��<�h�BB�U�jh��'@���щ� &˔`�'�� K����	�'����'�ŝ)�4a �gY�D����'�(���k�Y��ÁB�$1�
�'T�惃��`�ˀ1Jz9q�'!.�aHz+�a:�"�'�M"�)��<9������h^�������4B�ȓ*��x�#'U&E@ĉ�M��BI�-����s�`�/�" \��)
�;+�вtL#�K���O0��u�֎Le�z���<\�=��'R��" �� �|� �(�%.z<��'��%h*�j�Z�qѦܦ���+�'r�Xt�P!g����(��}�)�'!�è�Ra�v"� X�S�'�$�r�b��TI,hs�d_:S$���'j��p��>�����+�K0d�X�O����S�O��9#吮�f��B�k���0�'�$��Oɯ"4�,4/��0���(	�'� 8��럝 �j<��Y�Y�I(�'�h�˔���-;3 F�)4��'�Fya�C��p)P���I� CTI
�'�< ��Unu��"�
 q��=��'IHjR� �"���K�dT
01�y��)�ӊm��5X�
F�c"H5�bF�6O�C�	!o62���ڎ�ZLBת��X8vC�	��K�Y�F|��J6ZBC�w�R�s$�E�h`p�5#ɫ	�B��		���	Ӑ��)J�dQ���C�I�rq��a&4!�� ���b�(B�I۟0��g&�&yY��� 
ڎ��!,��hO�S�$�U��M�4�:|�S�Ȅk�B�I�K�|���C��������PpC�I�C89xQ�½��mAUXC�	h��1�@��X�ZE�ь2�2C�	�s��h�'�+n�� O����IH��He@^�vf��۶LD9_��1ס8�O2��O"��$X%��iG�+C+�U��"O �S�4���吡a�T�s1"ON8�#)B.<Q�c�eS	w
�x#T"O�襮P�[M��`#偐�PD�"O@� �DC%��qkSC�i�Ȅ1 @+�S��y@��fp��B� �Ui�yr�/m_�@eD氁e�٘�y��I�{���V@�; �I�J�&��$�O����Ɋ1�
�Y?M��	@h�-�!�$�<�$Mƭ��_�h��["�!�n�D����6-� ���	��>�!�<^��D�r�G�A���S6թo��	V���Th���[�u{8�k ,��'gƉ�'�Y�� ]%l"܄��g�0����'d�[pi����Y�iKXĔ8�'��p���O�f(�Ə������׌�N���b�'~�����$p�����|m���'��kw
+6�2mQ&��s��,��'��	U�)���%A2G҅MA2 �#����[��c�(�w��l�!bԋT}����S�?  ��ԁX��A���#�8�a$"Ol�`��V����PCX�B��d�����	�d�j0a��I�Vx�	\�3dC䉜>֦�2$O�R�$�P�e2C�ZDf&�7R��i����$Օ'�ɧ���D��^!j-{'I�(R����v�_ $!�D���A�-�bqТ�I9`!�5?T�aa2�E�T{�- "*�{�!�R@<�v�A�i@��d�Z�J1O.����P���0#�^��R��(�!�d; ��Q ��Y,$f}��J�@!��Q�V	x3S�V0i�4S	�M!�L���A���
��x�%�#�!��'dF��'I?�XH�G��!�$O��3��g�0�r�ʯ8V!򄀽?:޼��h�r0�'C{U!��ڡb��m`G��":Z"$J���i�!�d�<����dE�X��ĳ����!�䏗G��³�S�<K��C:E�!�ę�7��q.ԣ\u)5K�7�!�E-�2��-Ңj��;�DF�B!�����DXUK�*���@3�!D�=E��'�^����V��E��!�+��'̱���B��i1�Ӽ%��Q*
�'��cv�+w����1���35��
�'���#��Y��1Q���>)�"�z�'�n�*��:1Zqz�"Z0�:���'�m�旔Xf���!�$<+�'��$k���k�4~[L���D(<O�he�V�u���fk��5���C�"Oz�)a��%FB�m�C�G�d�E�v"O�A�`���C�~���@'W�xz5"Oɂ��>3���CD҃Mv�`P"O�t�ō���T�F+O�Nm�"��I�tG�B̹;~R��cśPh8=������0=����r�`���+d�ּ���S�>3��<9�@�`%3dIҵmq��h���l��Gx��)b1�G|�P����(���a S{�<���9E�V�ADՇU� �JM�<qedV4���Ę�%c��N�H�<��d3t	.��dN�#)\%�C�<	 ��uN� �ԅ0?���XԤ�I������%�4 ���8$(�c�Ո(mD��S$?��E���2��5N�t�JԎ>�^���G^0��OZUj�HC�^X���<��A��M�!~�p9�FdD����YD�y�Ub��N�D+�']��ȓ"�Tm#6j�״v��0Y�ȓKE*��FY6����0l܈9"Ȝ���H�I^y��Ov��ْ׆���&q�Ι��y�K�]���0��1��*�Ⱥ�yR�E���1�N�{����$��y"�Λ9+��#$��n.r)���Գ�y� {`H�cD�'d��R�a�#�y�MF$��)�UƻZ޼��F7�y��|�T�lD{�̆�;��C`Z�U�th9!��"4�ўb>�&���3 L�Fz1ҳ��-�F kG�>D��8�M�B��]��M�<�J�Xt�0D�p�e��gcT�F���/D� 2e��# w�)���ӌ)�|E���2D��Jƥ߆7K�(��a�.F*��"%D���wA~
��+�P��r��@���)%�I7Q�V��RcϨ���4
��[�C�Ia7 E�p�T�v���ޕ��C�)� d���H �Ё��=wh܋'"O֠Xe'�1_��ٰe�T 7j�]cb"O��t���sU�0�$ۀz�l�V"On����E����C�:/�
P�"O�ɡÆ��A�h�JD @0�$2��$�Of⟔&������7İ��7i��p�bl4D��" Ԙ@�f�ˆx7:uȣ�1D�XX��T6cq~��+�&(�8a�V�)D��� (@��$��(cbx w�&D��P��]�E�4@�:Kn �� �#D���A��=7P*�K�0Ohج��F"D���̖�9�$E��B��+���9�a�\�'�r��iK�w/�yY�*7u��Q� ʇ*K�!�]���t'�V�P\#⨞/<�!�$�cs�=a2��0ذ!Ņ��\�!�P�"N�w	����dM� �!�D�&`0ġ
�h9f��Ԃ7��@�!�d�#��C��[�M���d�%g�!��n�^��g��w�"��u�/&�!���$Q���8n��<X4�V�!��		Pe �Z�A� XR�H��m!�$_8�a�b�F�|�t�;wH�{g!�d��`	��Gb��b���*n�/D!�dځuV	R#�Z��Q���B�*!򄛉T��8��%�E� ��K�!�D�X�ʹ)Jo�}"�b�-OD��O����O1�1Ois4���l�� � �b��"Ov�;�BO=�����A\P�ŉ�"O��)�����BU�^�&d�U+@%�S��y2jô*��U1��A�~�@����yB`5#/��v�£^4�'A��yBg' ���C�˅4_l!s��U/�y���)+�L(�.#�Q!0Ę$^ �'��)�3扇:�
��R�F `s��icLC�I O_����!��>��!��23�"C�ɣ8�������N"~A�BV�q��If�S��y��E�qeF5��eM�W��� �Z��y��%S��i��؊:�U��۞�yr�G-H���P��R3�~WA��u�ȓ0#�4��X�r��h�N�>��Fx�|r���Xn�$[��3�� &�1P�!�$�x��Q!�����LAkF��+Eg!��%�����8� � ��d�5�S�O�V�{�s�Q�#�OS�c	�'Y�h����vX|��nܪ|)�<��'���
򁍥{{�q��h�$9`�'�@`h�
-]�L�+��?c�$�h��6�5��[�h���Ȑ�d�i�K���B�Ɂ-8�p��2�����Bs�b����e�S�'��	�NI2W��G���ꥆȓZ'� �@��>?��@��V6�tE�ȓ;L�i	TeЏb��ٳRKR���5�ȓ�F�"��I�L���8~����w!4p
f���lZ��c��<��]E|�'��>uPpW�4�n-;�ϹJ[BA3s+%D��������%��3=�dE�-�Qy��S;:��5���Ќ
Q�8��LM%aD�B��?[��CC�^!ba�x*��V$t�jC�	/3D�q+3�Pl��d��Cڹ
X�C��C����2ᕟD��x�F�!#hdC䉯'H�d
�&D�yG�T)*�
C�ɹvv@�E@cA��U+u;6C��r&�����,O�����Β
tc�4���XF���V'�RUʑ���*�k��-�y
� i��䀷.�����B�9v�*�*O�-����T� ܉������#�'�4����m_zp��/@�K�'8�`�8JD����L�(;S�U��'�b��!��v߄b�-��3��	�'|�E9��p��٘Wi�La��'��T��*Ӡv��\"``�*�JY��'�t�'���P�$�IGETX&���'aL�'�PQ�,{��]P�R���'b\He����S��_-y�V��
�'r���Q�Y�R]�k��t�Ȥ�
�'r�2�j���j���rf�S�'iX|�W��\�@#��T*��T�
�'8p�FŞ��E@���5�(�
�'^�D��d�.jp:$����z�:��	�'�z]3¬�1[,�"G
���2	�'�,`Ȱ�Z$x�ڠ'"�*!��'�X��q���Цe[6�[����'��aK��T�)3th�4�U�R��%P�'!�z��_F\a�4�8I�����'��ည�=K@ԙD�ƒGd�$
�'����ӟ&�)�B�Ͳj��]!	�'�+ �C����Bb�h갠��'u�)!����x��m�.,K�x��'�\��
M2X��ݓ��G�lX{	�'-��t.]\�>�s�cE��@��'�<�[RK���y�CŃ��	�'xx8�læ
�CEF�?�����'�I���#R��sA�s�z ��'�plx�(�}bA1�撌c?�%H�'*��$��yN�IT �)U�A��'ehq)F�ʶ%n�@��7A:Ec�';����%]�@ԦH�2ϐɻ�'� 
�Ν�8*.m
d�Y"&�f�I�'����FE�n�6����[)�y�b ����O+��1P�L��y����3�nZ�d��B��'���y�#�+?Z������PYj�؛�yB�؁t�$`5dF?�4q��I��y2c{Z"������,œ& ���y�
4�҄�ޡ�d�+U�ز�y"���|7P41�đ//�E#�y2� �f*�ՁG��3َ�����yr��|٠<9��p6��ܺ�ylYD4��`H�vVB�:�'W�y2!ŋT4�!`��- }�t�7jզ�y��f -�f��B��y:�ɏ�y�����@�E�Q�:q�mۡ�W�xb�'��l3��B$lQ��E~�L
�'иX��OR'{>�a2FU	{�y+�',��2��'5���C<c�$	b�'����ߖP�V�BJ 8j�  Q�'sx��1�	k�$��r�[at�	:
�'r��IG����(��<�TK	�'E((#���z��En�$_R�Qb�'>n�
����*���2�&�,��4��O�q�ۅ~�D�;�ȻK�n	� "O`PƎQ3N�UA��-z8��YA*O^Щt)		��(k&l��=�HҊy�_��	w�O�J���U�1�,s�X�.�!�
�'�~�c�i��{犌'���'��и���S{&� �-��>D;�'Б�,!���#AҶ@βP�
�'�<���_�c+V��/�?m|hq
��� h�#���,P|蓦�1m���g"O>Ѳ C�{t�ړEN5u>�$B�d�O����Oj�}B��)�B=�5l�kgLT�w�\�<���;�h��M<�X�X��DD�<��B�P���!���6�0�o�C�<�ٚ:X��Qnȏ̊�B)�A�<�������vB	q�zd/�f�<�S�Ѯi�z�
'��Q2s�]}�<A��޹�ܲ�� y/��A��c�' �I]�OژI�5�I�P�0��vK���Ҩ�'�^�G	P:�bi+��M�2)�9J�'�x�.Ԙ8Z=�������'"�m�d	�Z�\���'96�=��'���J7�K�P~x�x�.@:��8�'����%�J�#�(�����9����'�v aЁ�j�<a�B�`���ˋy��)��R�vM�͝}2�Dc@�P5��B�
/���!L��|�UNN�~��B�I:1˪�τ�"����&N�i�">!��	X�i$j1 q#�"g�"�J�K`�!�dn�d����4�i�$��f!�d�4S��� J�R��0¦-� KZ!���Jt���r%O�S�����f��;=!�$�7�y�%
�F��EJ2�ĘVSȣ=E��'b`��$��@�����c��4�
�'M��	P��<U��XĤ,J��� ��$�OB�d3�'8N�a��8w��]ZEGB�!�|��QR��c��U��XZ@�_ ,�D��ȓR����0*�H04�kN�V�
��F9�]��CZ:n B�T�(�D؇ȓG�:xqFhΰj�6���$T��ˏ�����84@��dK�a !8����q-�B��-YP0rvh��#~ �C�� ^B�pA���C�ݺ, ������USFB�I�A�@�����ky��b�3|zB�I<��&J�77�%-4NB�I5��ŢV�f`~%���V#Y�.B�#e$V0�e�١ �����O-({��?�S���� ~D� �  �oJhxv��	i�!��I���s��F4Q��P��!�\���<�o �]K|���d�!�$�>D���
!V������	7�!���=:��
AD�E��L	�W2q�!��\�E���J�ڝ�ʵ箂5{!��!��e��J"B�T��Oag!�K2ED���v�I�)� yZ�^< �'|���h�q*��S�CKL��,��'}P�r��5�<=P���!A)� 1�'�Py�� [�a�H�0KN:Ɖ��'�$�C���O�HYX5oߗ]����|��4��'8��� D�: ����k��ER5 �I�{�6Z����I_�ɗh'�4��S/I	��ئGW>7��C�8[z�ţa��	Mz�;�-W�8��C�I&J ��Ie�O�bu���S�dC䉍xS ,��"�l�ұdU�BdC�ɴdɹ��U�x���ba	�d4C�I�4��0�G��m�OE{�C䉒z1�q��
B�V#����D+)�B�I�P>��G��Bo�9��aB8�C�ɖY?�ȁq�ώ��M�c#�f��B䉭Ԩ�05�D'r���C��h�`C�I�M��Q˂�DPAaǥd�!��=�Z��G*T-b�$� G@v!�� ��ȰD�"�С�e��?Sm^h�T"O��x�#/�d�L�S�MZ5"O��c�!��(�wj4O�P*D"O1�ca��/}y�gjK��@�4"O $)�T+� �EH?"!�� "O�9&�9`�q�7�J���j�"O�$K�ĉ@R\Aǂ٨� հS"O�\1���!lr,m�g�U	F�Fa*"O,��B��Z'�e8pό"�����"OL� G>��b�C/S+j铕"O*0@#/�4^!��~�"�	3"OT����	 s��2l5�8�s�"Ob�9�)հlp���+@�?��!R�"Ob�K6��VQz4��Ʀ�\D0"O*(ʤ+V�R6�Lkb@ԟSހ�y�"O��	�FY�D�n��РT _0�u��"O�����V�|8pS�D�{'$�?O���D�?bX�(d��?1N�̩�I.�!�d�/'��#�a/S��3W�3p�!�D�$~Y䔐� �p?r	��nI�3:!�$��Y�,�)f`9CG^ ��ڧW !�H�zp��Їj6R���.3a|�|2��h��s% Z�w��Ec�� �y���8��S �������D�yB�Q�b=��`Ė�ʈp*S#\\LC�:*�� f�F;�Ja��R&5��B�1�\�4#O.`)��J�t��B䉗�1�"�?�%iäT�m�B䉢X��z�.T�8��%��i@�C䉙.�R(��K��&�� ��Ѽ%H"<��] R�bJ��P�׀��F�LQ��E~\�&��s(L�
I�H�T���H���o��,�B�GJC�P�ڙ��1ؘ)�+�����Wg]�fFvd�ȓMPⱮ��wFԘ�i���m�ȓ�@ղΑ�(x�gǋ%��̅��\y��uU	Y��Km�m�Gh�\F���Ɠ�XQr�I��N�̈0������ń�I�L+�h���P@���P*e�ȓg H�I�ڌ]tؓ"E:_������ٺ�
J�hq<������VȆ�{[2���f��3+�K�]�?�j��1�*�CJ�+����#k��-N��ȓ#&���a�V�d"K/�:�b�"�)���E5W'����p��m@6�i�<w��=z(�]"a�@���XX���`�<�FX"Iz�)�!�=	�f ����`�<Y ��?kư�����t��v��x�<���+� �S�NWunTۀ��o�<�H�$8|��`2^ҥ���j�<!��Ӱ$t�[r�ŗ�f�Jc��<)+Oh��d\]���Y͎Q��Hþ_*!򤗎@K���ռ1شiWI�
l!��w. 	���ߖ'u`���N�g�!�䈋L�T@�J�'A=���D0�!�D��W���6jʢ=Ƭ5�F�Śl�!�d	�A�����"�L�$�M;i�!�B}/H�s�œ"٤��C��!�T3iN���莟uج	�̂�!�dI��謂(�\����	C"!�\�N�ze"��
x����� !��(^�����< �L��!�$�~��H��I�4���`!�5\!� "6L�Y4N�|��v�R+?!�� �uk��0}a���o�o��H���g�Oaz}
�0���q��c�2�k�O��5|O9���Q-G�UcQ=Y�,A!"O�{�lj"����k� 2ip�"Or)��"N\���PTA7RR�1C"O:ĳ@K���Hz��E�M�6i�!"OZ���@HPf໖l�^�~Q�"O��Je�G;H ��fZB�ve+b������\�ON>U���؛U�} 6@@= , Q�yr�'�z�A�^	��)E!��_�f�b�'6��U�D������_���#�'�����	�~d�u
ѫZ� �'�����ډގ��я��L����'���U,�:�9P�d�C����'6h}ۤǒf�~U��J��,���
Ó�hO�1㒠��FCD!zR
M=_�<j4�'��	�2t14M1W)��z��YE��C�I69�>%wb�	���D�W�m��B�	+#ɰ�C�CVaΞ}2#�Ǽ��B�I�imܱyP�	`	�Î[�X��B�ɄNξ�z%nQ�d�F]�pJ�%�C�	��2W`�^��]�o�p��C�ɤ�Xy��ӝm��q�ե�6C7h��$�O��O��v`�:{؍�m�`�X��!"O�42�m
�ci�Č�=^@	ʅ"O�\i��@=xj���S�X�����"O^\���F4��*F�s��e�"OF�(���.}�HЛ�ǌ;d�m�3"O���f�f�����3L`p!�"O�dHĈ��"-I�^>t*d��'���|��O�A�@ �MW�|x<!: ��%�yR�S[r����$@xά�"�y�ʐ=W�����J[�j�j��f ��y�O�Z�pQ�dNߜY�E�8�y­W�5Xn�RtlK��`)% ��y��^x�is�&ݧ*� %LN��yR��>G�Dd��A$��1�$�,�y�	+j+|��6đ�7|�1Q���y2.ݱ?
�qRa>�]�C'��y� 
��~IQ�7
��m�bh5�y"( A�<�֎
�0�8S7JK��y�*@��$�BC;u\HEI5�y�C�W������/s�b��A���y�C�3(y�ժ�k`b8�V�3�yDP�dR�@"�,M�f����
�'�y£�+)�B��¦<f��[��ñ�yRL�&�`賂�=]d�,!���y���Y��Ҫ͍�����.[��yb��E\:܂uj^�kq��*"K�%�y2���D��ӏlԸ�P����yb�y��j򎟣�q#͂6�yr��=6�����C��	�^8�jL��yB �GYT�d˥} ��&!�y�GШY��T���s}��ڂg�9�y�l�08��m'�T�?<h�%*��yR�;C��nA7+Y~��Ԯ�&�y2l�y�Ya*Ǎ0YDk��y�'�w��Q f^�*H�[�G^�y2B��e=���g˟r�\lYD%���yr�t��q#�	��p��ӍM��yB��,��q�P���x����Z:�y�b�4a�
.�ڽ�I��y��5Kq�$+e	~�F^��1�'� ��@T�����giգ6�vU���� ��FN:�t{g@V��"O�	��bǖ�T�*���,-�!��"O���W��Gո�ŀ�?3���"O��N"Ȁ�銏w��ѡu"Oy�&�R997��.��b���""O���E�:�"�*N,�Z��q"O���g��Q?8�ۀlN�I�*M�!"ODAP$D�q�%��E=l��A"O,��-�XdJ��LqR�|�U"O�I)�ӪXWr��w.̭k�*,��"OԼ�����5����'��0�p"O�\���C ]��E g��%��1�"Oz ���,ĸ���F�c䌸�q"O�</��,IJ1�t��/'LlS�"O̼SfJ�8'F��j�)Qz}|�"OdX���i�ۓ�� -���"Oj
�6F%�  ΄z@�!�"O���)���p"H�0`Ь�"Ob4s'#��.o�@h�稞�O�����PF`�ႇTְ����ӍK�L��#2��j�US��˓
ьE��Vp����X{�b�F���n����l��0�/}��P�B/R�%�E��K��p�t/F�h��4Yp�;g$ L�ȓlI��s�e�- y�|���ʵT�܆ȓ:�ܰ���?N�Rҩ
�ļ!�����$���\$�se��Ն�d�֩��O8iMT��� �n��Q�ȓa؜9�B�0Dj���@�%�����9����+����r���F�ȓ4�:�2�CD"RF���e<E�^9��/B.$��`W!,�089��DB"��j�Lً��	�z=�6GEʀD�ȓZb�M;.<2&L��	߉��~f�Z֊@
=�J(���\�0���-��������"ܬp ��HǨ̄�p����a떭NΨ}����±�ȓG���7c�B)�3N�'�<��d�@�1�S;������;�H�ȓ?p�*�cߍ=�.ej"�&$�ȓ^v������������y]L�ȓ�Rc˄�ma�eZ�߾r����ȓll散��J.�b�OE�FqD��ȓr�
����<n��E�[�G-���}�x�rDM��t"���?��h�ȓ���T��Z�q�O� 8=U�ȓ,�P���B�&.��|QӊH Ojp��ȓ?c,�� ���_$�`�"�FC����&����IB�6mha����%n?.%��H[X� �!Y���(��_*���ȓ/�V��w�%%�Ͱ�N� ����r���CF����JA�� ��ȓ;��O2�pc���(5�<A��E�<bl[?^V�pP���v^XI$G�j�<)�a���q��`�#}�>��W'�e�<y���~i�ra��"F@ E�H�<�>�� @T�u{ơ
�#n�<y!e�4:<wd��t�N�� C�f�<锣�
��9�$d$jQ���w�<	2G�ż�8#��q L0R�j�<qS�D�C0�#�����^q���^�<�4j�mߎt�i��UpB����B�<y���Ps`/&EY��C�"�V�<�cT!y��q�$�h�rZQ�<� �qj�
�0�ZD���ڮ%`��@�"O��% ?]ȥ��,��Gp���"O�9��D	�\K�	W2p�˗"O�J�jqԾ5��(/!��S"O�a����g�~��HJ$N&���"O�j�A�>�I���c	��x!"OPh�A��� �!��[ w��-sQ"O�)����61�@�Y�S�ݪC"OL\�ͪ^d����A��O��M8S"O\�	�I9B�1�d�n��"O��ƥG1xK�����z�|\%"O�}!�ꕠcM����2��!��"O5e#��K/��+�4`��Lٴ"OveDD��c��$hr+�d�I+�"O4@�5L�3H:�}�1̊7���"O^u���_�,��MɆ���|i�"O<���SwnX��T	\�T�����"O���Oīqv�iw�[ ,��:�"OBCģ7}̙#1'�GDs"O����_y�I�Ǐ�t��dY�"O��Z���1	��U�fV;J�L�"O�i3F[7Wo��"����*�bU"O6��S*���$0)BDʣM����"O8)E�'Ĕ��BDK��8#�"O�yZѪM ��� ��fes"O����TA&�u��L,/>Px2�"O�X���ɮ\P����F7lqZ%"O�Ⰵ�%w��(��1��Jt"O4�&��q�8+�d�����'"O��S��=;�L`�2D� 7E��""O<h�##CK{"��G�]\*��"O^i�g��
ܕ�p$�3ǦYH�"O(��:{�dJ$G��
#J08�B�	Ui���s��dl�Ĉ��G
`�(C�	.�-1�J_�|6�q�`G:-�
C�ɼn��X"F
gf���Ŗj��C�	7j���a�J�֐�z �
�C�i�%N�4U}�����1�LT��o7D��D�v�sD��De�/D��c�Zt� P�V0��
0D�đ.�?{s�d�����;�O/D��S�m,��M�H�'#��A�:D�C���$S&��;m
s�aPVJ:D�(��C�/OU��u�S��,�7�7D�H�HPv�Z<�6$�_~��
w-5D���1Eل �DU �7OR� sC�8D�T���W?�!���-}zt۳�!D�0k��GK�ȣF�㦀�2m3D���/��|�H�tEU5(f�c�;D����V�dH��Q:qR#'<D�|�1�ݖ$_�+E��)]w����;D�(���8'�*AB$(�����8D����It.2DA '�1�F��A�7D�L;��� Yk��B�	ݬ� `��:D�и���&�G�"t@�a�O+D�(�#�W�r@��.�3|pP#�*D���� ο#��t�+[EZ\Ҵ�(D�Ђ� ��-��,�te¡E+�10��&D�|y�"\�v��@L_+Q����!$D�����&Ҁ�觅]�1��!D�,p��ȣ8n� �hڭG�|A�r�"D���c�*=�%�f*Y�!'T�Y!D�l˱j�+��s�/�;w1~x��>D�D�Ǝ�B�uA�! �S� ���=D�� 0���=�7�J��ݙ�"OV�4EC�J��	�cP<3��4#�"O���k8r�ʱ�Ͱ:�N4��"O23S+5<��� ��9�"O �*/K�k'�a�3o :]�Zd�"O^� ��3�:���An�p�"O�����l^Pp!�E4X� 9�"On�ӴC�6C;e�Al�3;b�I�"OJ}(�e1h��PhS(IѸP��"O<�:�ҟ[VB�q&�R�(�x&"Oz��ӊ�?Ja6ͫ�c�	\�~ �"O>� %�y�"u�ƉUP��f"O�Mȑ��
�xX��R���JG�'D�t��/ё
� �äh�P	:!
$D�; �E;;<�<J�CKK\95">D�� ��N?y	N��v#�:m�%4"D�0�(E�E�x؃7�m���k�!!D��	��I�B�Ļ���\xz}j �$D�x+���7w�PP�H��{|4����>D��0���U# �x���U���I�=D��R��.�09�U�sֽk'�;D�Ъ@H��"��р�,��$2� :D�hr�j�1a���I?߰d�1F+D����kL5h$�F=1?�,��e5D�p�E)F&@/����A
r���1D���T	Z9���Ғ��%y�Fl�p	,D�[�J�*��I��Fq��?D��q�*�5;��Q�퓘'l&� u�=D��ʒ��[��@��葓)�����(=D���w�K�K$ܝ���~T�?D��k%����=��.�k�T�=D�a�mӝ9�pU�Vn
n���1Vg6D���v�5��I�&S	w���l�<	]����n� n�t��5fU�i����'�0Q���<zY�C�U<��y���0A� &4-20H��0��ȓn��7Ɯ�B�$����MHV��'�Ak0�UhH�P�%_x�¹��'�b芢�
(L����2[�Cp���'�q�U���R0��D�A�G�ȅH�'eN|�sj֣x+scm�L�j�'�%�j4ci2�#Äߟ]���'�r�	��8/�� ��'���2qx�'^����!��,ݴ���ǬU���' ���Ƭ�l�����/A9���'Vʹ�p�ͪs����!	L������'F��4@��̌9�N��ղ�'A�=�.N�w�0t���/
�����'�}0��ǃr �p)י+��U��'�U���6 �ԑ`�^��j)��'�f�5KCy��4�	��D��'�-��*L�x��y3m�+���*�'�~�b��"<�`Tc)��8Y�'j��{¦�W�L=�D\~�8u��'X<�QfȓH�а;�Evx2�'.V���k��j�X��ᔠ��'��kA�Q�$�Z�``��Y�6*�'��c`��Q���a�E�LQfЛ�'��6��,2̆1��݋��Q��"O �dh��L�h�Xt	�Y�iT"OX���́�w�(��'EaIDbv"O�8ɢl])�"�3��-4�0a"O����N =:�Tzf6->�J�"Op	�t-�.���xd��	���K�"O� T�C�P�NK�x����G��)��"O�����ʟ|���4
@):�nq�E"O2�:g���T��5��i] wjX�"O�p{0��m.v-��i)fLyp�"O���ZL+�%[�JKEz�|K�"O(yst%�/w`Ċc���'I.���"O�i���Y�jx~�����9C��a"O� Ӄ�f	|��F0
A4X�!"O"1��ʞ8+�a�ƆD2|���'���M�|XSG����'b�����f�<y2���|�t�b�'WL����X��1� �CNb-I�'�ڵrAݭ^gB��2�*�,ܨ�'v6�A$�4E=��"���)�HJ
�'������O(.ݾi�I�%>��	�'ņx�C�.8$�D�׊��P�
�'�]8��ʊ�GQ�E���I�"O6�sA��*7��=k�����H�"O��0��A��84��T�SR"O(0�`
� ml���0	��I�"O�� d���-|�U	�ʄ�`(��&"O��§
�7N�܉�	� O��s"Ot���)U�[q��GS�R���"O���τ]R� �7��P��Må"OR�����!G 1{'&�s�H�`"OФ
f��=�h�2�啍U�Q��"O�l���_�^�@��ߴ��1 �"O��C�mC'm�,��٘�ީJC"Of�Q�fN�(���nD!��l"O�y��BH>H�N��h�F"O֔��c,��̈�=�Dt�"O�6˒�/�x*�%C� �|��V"O��0�R�.`$!A�[@o�H�"O@�֎�x����8j>�"O>��u��(��Ԡb� ug*쀗"O>es7kP�DPj�C�m��?���C"O� �R��\e`	��Jd����7D�Tӡ��/(
���ZS���%f4D���Sg�2i��go�#%� �3D���g�=X�@�`�D�]�U��(1D��2�aѿ"�IY �ވ��!��&1D��S�,Ɩ*�@P��	^�`���A�/D����݁5�,ܰ��ȍ,�� ��.D�dK�?�,���;�
т�-:D����V����wN?|j�0�7D��b-�qyN��aĭ!��m9D�lx���
�-�e8(!��<D�@�7E+UȌ+7f�"p(�2F6D�@p�R�����"��$6��$�4D�4&'[�%��W+R� ji2D��{���z���f�� o��2Z!��<�N��5��%r0����*/R!��I�l[�e�qK� �C�W.\7!��2�yE`�6-.�`pDZ�H�!�dQ+m��w"S�WA���˄m!��޸Hj�<�b�)Z�>�A�'9E!������zG�/��j&��
gZ!�d?b��J���� �R�Mڕ@L!�D� c+�ѣ�k:joz��v��#0�!�䎙Cn���NF�C}�$	��W<�!�KoP��¤X5[*lR�,X&z�!�ą 0��tㅪos���!�4@#!�dL�E`v%�e%�p�M0!�%N
!�d���IAd�׸V��G	U�_�!�� b�[7�ǆcڎ�3���V�ʠ	P"O`�S�Wz�90����s �:#"O�Xj
0.@���0��o��yxf"O�M�#+E45� EX�E����"OlDCr �$�4Ep�M׋4]"��"O�9�fa�?,V&�q��x����%"O�ݹ���� Nʼ��Oߎk��[ "O��"��8�=��@��N�"O�(asA [�|��.b�d��"O�@��0��{�M�<��H�"Oj$zc۶&��5k�M_ ��MZ#"O�5�P,�&����t[�\לi"�"O�Ð�?]`ˠ��f�� B3"O�X��N�8\���ƪT���9t"O(���S�;Ę�3���	���"O�屁BX����"�V4f�^萐"O����Ȣu�*��3HE��A�"O�ᤦ��E�� �IZ#?����u"Or�AC�&_�RD:�IOnPa�"O"$g�F��R�rv��"O����a��Zd��qi ���"O:�"��#}�e�pGW,BaB��D"OD)���� WՒ�(�/��t[>��"O88���2dK ���@������"OD�{s��qe�����l;���"O�Q�  )-2����1
���"O�ȁ&�7Mq�Q[�ꏻ[8��P"O���3��=?∙���P�!jʑ�"O�|���ݹ;yb���Y�[���"O���"ဃjb (�)ׄW¤�"O�!�2��&� @���N�
b�� �"O�a�U����j�aG�V"O��R+S�Y���F�S[$���"O>�jC��#d�rp�d��rV��d"O�%��r�Pա�&����H�<)Q��A�6�Õ��4-��� �BB�<Q��q+.����P6t�(�@��Jf�<Ѵ����h�*���b�끫Fi�<	��P>�:|��A�V�@�E�c�< &�.�d���p����.�yR`׀U^h��w(H=�������y�Ok��0S@+[�7��M��Ȁ�y2�B��f�C!c� w���y���xv.q��0 ~��v��.�y�*�,L%(qIRi#+��҆��y����w�)k'�	�.�t	ۤ��?�y�ɁW��t�/�DaTH]>�y��)TBd�)��F�=t-J��y���F.|��,q&��4�.�y��C/gD�$fݝ9�@8T�ڟ�yr�܄Q�$j4F	�7��)y��H�y"F�u���DB92�(�	�"���y�-ڊ=�Р�`�&�z��T��.�y��G�v�:���-� *���K�G�y�Er���O�r��<�cE[��y��'P��	p�΂hhԥ�� @)�yr�';SL���4[�0�Aԩ'�y�d�_�Ȑ���	UO.�)�`���yr�K�e�<I�����\�lu�����y�^X]j��G0R�v�H $I�yR�&e���8���H5��J���y�L� ���Ĭ�q�`�	cE��y���1R�~�P�&_(�hػ���0�y���%u㜁�QNٮ��$Ӕ�L�y
� ���h	H8���y����"O2�Bێ�[Up���l&��e�3"Ox�wF֞r���C\	;�0q���L�<q��؁y)�P�%2<h�e��S�<��I�6hݐQ��=1���ѣ�Q�<��lK�@��,σZ�r9b�ɘW�<�6��<�p0���'*;�ZKSO�<ɁG�^�^���:g���Zf��P�<9�]bQ�%xq��n��y�FDs�<�t�1HU�z�h�%T����p�<��+�z@��jr*��'�.����
k�<)�Zd��$���&�����P�<1��X�c�0����1Xo2(iA�GN�<��D�+T�.I��+�ـC�N�<ѱmIx�����:羭 aCQ�<�p
҉D]�HJ%kڃu��1��@M�<��BD$pj"N��fH-���EF�<�2Bݾۈ����&bp�95� C�<yU,[=d�v�qG�h�	��|�<�̍~��L����&o���Gw�<9���Q�x�'�[:�qDhr�<�d�ER����	-��`1
W�<�T�8�~� �h�P:@��!�U�<�TdU�;J,!E�N]�D�DI�Y�<a�.Ѱk�.�S5�؎-�� !�XY�<���\<�RIR6O��Ɯs��]�<�C�U����I5	��xJԪ@Y�<�FlD�'�	��J�m���:Wʙ@�<�#�.>�X3o3BB����Z@�<AaLؐ ����䉐�:�ذi �Ux�<�G^h�� p�ʃ�5��Y�bE^�<��`�z� 5y)Y��	 f�^�<�#��N�2�X��x��}ق�DZ�<qvdPi��<��C�,��t�Q�U�<a���:\�eBF�m:�i���O�<�A��Hv���Ĝg�(Y�	T�<����Ą�����f��I��!�R�<!�	�&���f�X�O��x�eaSN�<i5	ɥ�,���Jv����I�<u.��*L>[$$X2�f�ː��z�<���X�eH-QT�J�B��LC��s�<Qp� cĨ�g�j��)���p�<i�#�9B�dL2fh�X�>���[D�<ـ��|���qÆ� X���}�<	�O�#]����n��h�I0��O�<�W$=fy��`�Ɓ�a�l��!BN�<qw�ׇ}I�T���$5i�
F�YF�<AfD�ߤ̰�c\ ;��)B|�<і��5N��a�@��b@���a�\�<�ƥ�6@���	4�$A����f�[�<�d��]��ٰ��"w,�BרAP�<aC:�i�����BT��*f�<�uO¬v�~��u&�5���k�j�<�Qn��FĶ,a�h�Q4����
Qh�<Yte_�$<��ǀՈcv��gB�g�<!� @�Ob�T�7��	�r ��j^�<a��ܜ@4��bR�U�@C�PPE�UD�<9���u��T:�h�Z��!�Ӯ�w�<��hZ�$R �	V'ƨ����TFt�<��!9�s�܉Zh����l�<!��
�F�-J/S	U����n�<� ��&#V�@eG	7���!+c�<Q��E�/r@����x��3W��X�<	עڃjQ�-�*ۅz��;&fJ@�<� �������]	4)Q��A+z�Y��"O����$wl�Z�Y$>l̄k�"O~e#�Ӑs���ԡ�?$T!�7"O�����8U]D@���ذ�V"O��ۇ�ձ�8A��;�p(�c"O�b����KT�"`�/LҊ�� "O��P��Q]|��ף[�Eq|���H-D�0�b�Z�"���k��P�e�F�5D���FD�I"�� �o���%J)D��a�H�Y�L�{f�\[B�z
)D��8��!,����AKN�z:��.2D����n]�2hA��;7��ك@,D�Hc /v��x���Ǜa���t�>D�A��^�+��8+�#�v�Qj/D����+� x��[��F�(ڂ�`t�)D�\�V�L=n/�U�CAE�
t���`&D�8�P��"Fl`u/�	|m�}x��"D�\y�HP��j�@�Q�����.D��0�v��=��J�86�`�<I�(����Ui�K�;ap��
��E�<)H������������E�}�<�/%m��ڣ�O�49�5�Q�Ry�<�!ޞj�]��Ҫ��eK3�QJ�<a��!\y��(�?z]F<{�)D�<��o��:�����-L��f�[�<��d�3A
���%��!��p�<�&g{�����3����Jt�<�B%[�L!�-���m�^	�!-�q�<��[�O��#cD��*���+r#�l�<�A�1�h��7L�j�$�+ť�j�<	N�lu�u�5�։#�ёB��f�<I��L�w��E8T��Z��A���b�<i��E#�� �
��̠KF�G�<A� �[\J�ÑdV<)H�q`�\�<!B�Ҥ>4|�Bp���lxJ�Q�/�V�<�*\?`0�bu�,�����J�J�<��/�o�8�s�	I-R4�T	F��`�<11�HtZ(�X!�ގ^%A�(g<A��r�8����z!>5`�Yt
��ȓe������3���[A�R���I��
ZD��n�u��y0���xM�|$��D{���冡EJ
i��J�4�Uz�gY��yB)�2Rn�z�"�*�Ȅ��^���'�ў�O�,Y����*�4 Z��M��C�'�4ؠ��B?x"Er!b6g�(0*���<O*���nB1h�̠�b��p��"O�m�@�V �i�GK�B�$�i�Y��D|��d�4��)HGOYC��ɹ�
�]�!�$�GJ�pS��ҍM�f<�$���d�!�D��)+��z�M�\����O�!�dE�l/RIW+8 ��(1�k�/�$Gz��9O�͹7+�H��8Ԉ�����O�U����_]��1��:���f���t�$9�ӂ�$XY�!'lF4��I�~b�xI�:$��]"��0īD�߰>AJ���B#����P�m�\�Y���;�D,�S�''�!@��8
��Ѕ(!���?��#�S���l��9�3l�%r!H@�M t !��n�Z�gˇ}8%�G� X�!��߹<#����)ٴ%��q�f�Аk C㉺�z	S&/DH�Ѡh�~m�C�	���L�7g]=������^8gxC�	�}|X�7�M%=�y�C�? �B�	�~�4��7�F�nOz�Y�+S����TT�)�� ��Ʊ8b�$jsh�E��"OJQ
�Y�8?j@��g�-$����c��k��~���'p	��!ǲ)���B].Q���C�a>$��RC'�9lT�K�I˂A �e�d�-(t 㟰��	�wX4mS� ʆ"W���Ą�7-Z���4�$�'�ҽS1ȝ�\;(Ab7ND.�OΌ���TE�s�H��U�/�l(�U��䓪hOq�����[9^<�g��U��)�	d8��s�̝(Z�����}�#��)D��P���?Ph��>4�8���$D��3��0{��yj�k�B��,��"D���/6d 
q�S�+�4Tb��!D�h��F��h����<:��)  ����I˟l��Q�)�S'd/z ���� (AL� H&B��,��q��Y�1������2��6-%�LK����YɆ/̧e`�!�n+���'W1�x1��͗=8�}�6�M�_��-B�"OJ%)�TH����B�|x���Vc����'���s����`X�I��y#CƂG��4@-)O�=�cf̗>S~�*6��I��Rf�V��F8��8�쁶2ĨiX�k�I%�Q�G)D���Ɉ-�
%���7��V�0�V
OH����D5;?$�Z�IߚG2@����'��'^�����=.�T�ߎ_x I�'J6��u���bH��(� ���'P�0��$\ U�=����B��E��'B�a�O�OL��쑺7Y��N>��:w&I��G,*�(y�f�ӎ#�*��I�<Q#C
�A
���!.�2E݄xX�OX�<��O�7 p'a����h�IYI����O^h��bτ�vt �FI��)� Mp�'� U
P5Z\�����(Q��d2�F���*!���^B*:5�a�'��Ε}�<ٲ�eR5�N����Բ�!�U8(Ӭ�h��o�~D W U8S�!��2iV�:2����-��_$C�!�E� �T��3Ȟl�Th(���3�!�dK+8s�� ��2hР�P�d\�)�!�$��Z������-1Ą
 �!��4o�Z�H�V�s��5�$�ݏx}!���;_&|c��ϨH�J��A�t���>�CB]��r����(H���ِʒY��I��O�`�m�(:��$�
�`:���"O�"S��(����
E�R|n���퉰 ّ?]��?iƎ����K�,al8|O�aK<��ΐT`m�S����r1���A�<�㭋K�(Y�V�Ť4���8�gUq�<Y7���-.��B��~&i���Uo�<I"a ���@�蛒"0�H@3�]d�<��D��x����r�
d����i�^�<yB��T(���ć	c������V�<� Ҝ�pT9�
؈X�a�V�<�� G�]8J�;�ʂ�XD(Z��x�<q6-�o5"(�@�My/r�A�[�<��͎�%,�MKФ��U�p��[~�<���6��B��e����B�t%��{� ;L�qb�)d�X�. D�44�s��8Q����;����?D��p�ѥMF����,of�trį?D��yw@a&*u�a*L�D��P#8D�D肊�hu�� ��E:���:�rhYD�� ށ1�����(�u$��+	��y��\�AUPĒ�Dƒ}A�D@����1OX�~�G�}B2 ��c�^�����Iy�<� t4wg�,)M�,�����RbE��]�$���H�6r�G�2nȼ�ܧj���"OhM��,	��x�g�O��d{�>����' �O��@bB�/���
��W�x`14"O2(���=z�*��fQ�W��5�g�'�!�d��1TI	����7_�+�u��{rR���\�8�EM�>�^L�A��'Xf�H�� ��|�f�E�� Ʉ/��7��$GR�V���`��I	lp\�$B͍jC䉵>�0J�Fչ��$���yPXC��,�*��FF7>���;�=D��C�I�Js8�qD���� ��дl���r	�'�,�@�X">t16��	w~I���(OI���P�gq,ɘ��؎�ё�"OVUU,�_��	2�%�9�J�3�"O���%E�=5(d@�%�B/D�Ҕ��"O�m8$.ji�x�D� �҈�R�O�7� ?!/O1��=@q�Iq�&B_��R�o�3,;.C�	9U�Xp)��_�cZn�� ���'�a}��-,�){`����9�%��'�y��Q�J��dT��V\� D�¤�y�J*<���y��V9�j�H��P��yRÙ9pZ��G�h� ����yB��$H0f��0c��3��KQe���'�az�B��8��'�1@#����C� ��x�\��1O�*	u\�
B�"!�d���*�R�ɟ4��5�u�U$!�dC)T8f=RV`@">ڜh�����!��Y�b�#S��Z�h��5
�;�!�D��/T)qPeH�(�rd	a�O&�!�E�sW<�SAĚ�[����%$;�铽hO�h�X���#/� ���<��\�"ON����7Ym�$;҈����c�	P؞��uF�d�`fԸ6
��À 3D���S늷j%�DO�(��$�5�;D��Y��N:�]���͑W��U�g/D�����C}�uR��5l�)t�/D�8�Ԏ@�_����C�09���H4�.D�|��l�_!�2��8�-r��(D��;�����,�4� C�D8�C,D����a�E͚�S�-)&ԸL1�M<D�D�E�Dx;\�L��$��x���;D�D(P+Z�VNX8���8Q�H�F:D�1�䟵K?L�z!�A�=tmRf�2D�\�c���i�n_#Y`����2D��ӄ��Jl;4)� :P9��g1D��ɱ/A�9N�iȄ�Y<�&����-D�����!<�ht�V"��#�%D���!�B+$���$��%ĩ��"D��j6n@�07|�ӌ�?l�� �� D�d`�MN
g��SHC5k�x�a2d2D�l�u�������W2���<D��rFNŏr��[AY�x�� �
'D�@����7�^hQ�+uN\Ey0'D�ܱ�d�4I�JdAB��$� m�I%D��H k-������ly�Sh=D� ��#�h�`��%�
,<�L�*O���ED�TN`��s�??;z�P�"O�t�K�p[lڕ�;�Z���"O���mK���>&{� �G���y�%A	]���$/ܯ���:FCP:�y��ů_�x	۲��F�>�Qf@��y�FǊv��<����*=c������y�kEh�ȕ��%7:3�)v��*�y
� �0R�j˶k�Y�F��s�<X��"O�8q��DK�`���;'5� ��"OBip��36�����A`DH��h��@����\$@���3h،Ab��{f( a�V0S�!�ĉ*�x@��"�����SqN�!��m_�i���%���fg^$�!��F'̈́Q�����f���@ ݗe!�$�&5.�;����;,�V��JA!�aФ�0�R6���*5*V�"!�$_$}�z�Vl[?�>�8��k�!��2�D�r%���4���6�!�UpG��g�ʡzҘ��S4�!�D�%_��w)D	��`)�9w�!�$��E� ��'F\�~��0��D�~�!�䙴A�X� C�Ty�f��DlQ+>�!�5 1t�h��Y�"���2GJU%22!��9-�m��N��eC �@/C�!�䈄k�и��A�&p.HY�b�P�!�d��A���C[z�ء��l
 /�!����͒��m�>��p{��Jz�!�$ 8�ţ�R�C��(�f���-�!�d�z��Bv� ����seط\�!�G�e��|���	&r�� ��
�!�Q�h���D V/#;�E���Eu!��#�>�
�������)ă�z!�$�-_�n)C��82�R )�É6Dd!�d���0� ��$�7"ո�!��I?F(d3'��5�(�ඡ8!�Dˬhh�d�	�/��H�[?OP!��1��9��Ύ `+�,�@D!�_�(�*�� 2��r���~�!��M&�1r���9�H�4��7{�!�D�s�lLȗ��:�hx;mW�+!򄟐b\��8&#O�V�0ձ�̖!�d���'+������5�����"Onp�3�xY�H7a=�5�"O(��#E��-���W!J{�,8�"O�u1�a�Mz ����sh���S"O��Z���
���
EFo0��"O��J���EO -�&d�r��2b"O �s�M�^yd	�����P�rM�"O��KO%z�(�u�=�^��R"Oj�h�P���Hn/B���Ӕ"O&X�e	-D�ո'��tʳ"O�hg�]���Ը�+Լ�.)a�"O�`�v��}��] ��&�f,@�"O�t�G���%��f�%��عf"O��[��Es�z�r��2"O�-�����,� ��8,��� D��s�̨vup��d��>���S>D�L�`
3;U<i�B�:K�U�U?D���v�:A��C�/��|F�4t'=LO��ط��>"h��kAHu�1�ߒ[4`��k�Ԥ��>�Ü�l@��Hd���<'��X$GɌ��,�c� T����&'G�V�B|I$E�4?�\C�	wup�r�O��;�
��S��>{9�H'�G,��	k��� ��L<��e�#S^f��b��6%�X����]H<��Ț�5�h8��hz�F䙕,���
h �f�,���k����B/f�lȫӎZB�zȅ�I\����'�������4����x� #��%0��ȓ3�Z� �N�����5Ȝ(OLȥO>���+��V���&�k�O��M�G����RICf޿MА��'#4� ����X`9�+�K/�g��C?QTa��__�`�|�I9^[�hΓd;�d+C`B�P'���-��6х��e?�D� z��l�+l�8���+�j>l�3FF�j�Ƒ�VL��/����փ�=b�nȐ�,<�`�H���d��y;P��1Jnp��ɠ_
p�4Oڂg+�Eb��X�R �}9��״��́�#��?�h[����te��
\x�<�ĩI9(�S'=vxQ��1?����>|)�����f�89�倠{���������&�l����RD�%K�.]�w!�	�x�FL���M!�$�ge����,d�������~yZ���S�S��pQ0,m�I*��
{�`���}�<Ѣ��$�@
rʚ�j0T�d�R���A6�P�K�l�֣��M hEl�=°9�@i�.�v���I��	���K�� `F36�Us�lF 7�(�;����0<���g4��%!_��M�R����:��N sk����,=�t1���à�� �fO�*t*��#j�<�#�<§N��ɓ����;�Z�i�j�Yl5�O@�"���5��b�'����W�	D�k�Ra�D*�Ef�T�$�ׂ&JJl��'�<SG�'*�(aʟ��T鞭-��+#kP�P���	��Ҟ@��'���£�|���@+@7����$��ӡP�>��X�I71��"e��*h��q��	�7!v��Q�0�T��'J��.Obt�r��t#]��D��	
Q�G)7��O9��!Ǝ���	�%C�/� ؊�'��� �D߳���ggBS|v��`욈N�!K!�?tz:�H�'�
��O~���#�����NR�C�s&e��^
=@�E%��kG��DH�ٖ���?��b�����  t���oˎ��-�/��xۀ�L��OR5z1�	x
Q�u&ˋ.�*���'&�58�ך)(�|�Ы��Q�J,S�`�6`<��$�b�T��A�U �M3��/�O��K�px.��SD��s��L��>	�G=�
-��o0x���p�$rz���c�~B��6�'�7:�rM�f�Lx�<����. �5��1�\|e%�9Y����Y�SM�	{1�7T[�(�}2��*���^�Z5 ���KU�I��Ź7K��U���V��<�P�mh��PD䔙P�nP�f��M�޴���"3�U�N�?!THB�S|l%q�o�"�����*�r8�����>�h�'����G'��?��H�M�n�X��#7D��(%����Q���^9xR`h5?	��.B�z�*��0���.@�p�O�f�CA�55
xS��K� ��U�� ��A���F�9�Yp�� "�&$������ErW0�&���O��B�8h�)� ��l��a2�I�`�p�0Q�5���r��;�x5p�I�:�l�J�"O�X�0;
`r�.m
^H#S�i���A�@H��M�O?7-�:D.��w%B=�`�c��ӶR!�$ �Ԝ*��Q2Y�"={�F;�������֩7��yb"U��"���o.
�[׀	7��>��N�h�T�bBѵ������E��{l 2�C�IOpDM�ȿ�8�P��Q�4#=i��%>�>�8V��OL�PJO(�����&<���yG�B����#��yr�+2Ѥp#�`Ĕ��Q�����Mc�k����v�lòN� F��"}���ڴ�N�|栙�4�Ѓ;±��t�*��h�͖����9fX��i�OҜ,�.�`��+[(�k��Y�$DC�jjR��rk_'v�@��D�H7�hY��	7�bM��f�/
j8{��A��v��/}"(=me)��qAQ�~�{��<�;ǧ�A�zЂ����O�U!��'�?�d�\��h����|�BʄfU�=��	�5��!�"O����3�h2���l��$�a�d[>3Cj�0���h�^)�,K ��isG%tZ9r�"Ov��@a�cR
<90E�$�^��׋����A��C����Lu�شˡEQ�sU(�㰇� z�!�d�֚�v�(�9��ǉ�F6-��%r����
�=��=���,Ϥ�"e��5�]1�,�Z؞���B�0(!�qC��'#`l�gm�dv�)񇄊q\��
�'k*�J�F�7j?"e�w��m�l����c4�D���`P�C�,FUl����	0�C�I~�B!:�!��]��m֟�N1�i��bqO?�I�~��:'I�w��{����U��B䉳(:�(Q+�-���ض)�a}|<��#?��0>?Q>˓*�^�[F�E %%8ɰm��Zb,i��I�!��!A[���qCΘR�6!W���'@ƌ���5�1u�s�a}�%[_â0�"��4�^ ���\��'.�UK3�=,��і d0������7��ϧ�X�XAO��KCM!��0�����J�LK�L]�]	d�5�~����J5v_Q����bE�M���H�DCO~ʐN�ڼ� �A�%��1	�H����Kz�jbP"O�a���W�Uf��4 �7;������nvb=+E���N�Q��[/�q��ֲPj� �N��3wDla"�D�l0��ed LO�$)�"�0\�""@��u_>|�a��;Q*��f��a�q/6J��ge�ne�ą���:�!�S���Tm��dc���$-љ�pi	�!.���ٚO��Q@��u���'z�����e	�irUJ��y�%�.v�݉��E�TO��Q�U7MS���Y�R�su 9DA�t�@�,u�٥���9�j��P�
�o3���!��1�r�c�"Ov�qe��g#�x
dh��I���6���R���M&A���D�/jr�A�%�b+�h�{��- �d��cM̎@��L��N�0=��ǡIY(H[e�G�f!7�$�d�e��*M���B��u(6u�0��U�݁�D>\O� [���R� A��&%W��@S��+`t����'�&[����i�34�z�[H{��y��T/3����c��YG6zH��y�"��ѡ���6^il�5�A��!�wl\�{_�q�5�#_m�8��^�}���%?�`�wCP�� GF�� �X��`>D(�'��UU
�����	םP���v��t�@��0�,h�z�i���ħظ'$ ȁ�E2MH��"�+�A����N:�C���łU4V��Zth� 	�d�p�IY%H�q3e�(�p=����.Ir9a��NZ=J�)�Fe�'�"y��d�(?K|�`�F�W��=��f�(Y�1OӟN��PG��}��ȓzݴ�i�O�6�<�qI�2(�ɕ'���� l$%S؀�Vg6ov�<E�4�K�K0������� ��h<�yBOF��8��$�����KѮɲ0�j��p�8Nc�h_��43���yrbS��@��_�zs$�[�H�xb"�(�l���*K O�H���
��L���i�((���4�T(h��{�k�.�z F�^����g��p<��A�Jp�Ӄ&^!5o6扡	��"Wk�UR%ۗ��@9�C��eQPe��^�n �xP�E�|bÀ�0]�e�C�O�
��$�������!O��x�N���'qig�ɵ�>���ЊEH�,���P��'B�F�,O�l��,��K}V��Ӥ�Ux =�U"O�P�*@�z)��3���2y�ؙ1"OI�OF��`�?B�
�ٲ"O�J#��N.�l L�e���"O��2�$߃+�!cW�ٸVAF��"Oe� ���W���"D��73|	R"O��:h�:��]CW�T1 ]&X4"O����Z�5a�	�2�F7�:��"O��Q�&ʃ4�lEk1AR4��"O�B�,�2&�4)d�ù^�%�"O���I����kT�G���e"O45j�Τ.&@�����#�rT��"O��ԊM�W��=㑏�Y�H�{Q"OU@V�ߣTfx��苗gkR���"OԌ��b�'����7f	FX���"O��+#.ه<�\}���-��� "O�k��W�F�*G�3r�,Dy�"O�e�# �QӾ%)�b��)��U2�"O�E{���B삷a��=˔"O&|�T�l����$��\ "O��Ǭ�P����b�9d���B�I	Œ�ѵ�P:u�<�	2�ܒ(ՌB�I6_LN��a�ǽ ��d��CY0L��B��?:��cD�<+��x��2�fB�ɝz�z��oٴ<��ya�̕m�*B䉫Yň�7ᖨ\�JP��ߐ#}6B�	�d�z��!Aە�XxAN��+g<B䉪<�m��F�l�<��`c_�}�PC�	39���H�� u��H���+0C�I�4�XahҀ�	��EK�BW	c��C�ɐX��7��ad�)Q�3=<~B�	>M��PY����ɑ"�� E	B�Ƀz�&���4U�d`{�$��5(VC�I!9�I"�ڡL�~�Y֦��+(lC�)� n� ��S�
��'b�*0U<0D"O�c���{�N@��5FNP��3"O�5��Ұ:� ��/�O1�Ʌ"O���LǓG���xF,��v�\|z�"O�	��ŧ(&���A��7	���3�"Otx�%��>�X�(�����1��"O�5��*U*5�!dj΄%���!�"OF��C�gQ΄�p�o�8�"O��s�,�9fI���dL6 �щg"OZ��dϋf��g�B���@��"O~@����(3��#�ař�,2w"O5�	��b=+��Q�@�CP"O��!$��5k��L9k¢�"OF�� %�G�!�
R���=��"OpșC_�f����C<z�T�H"O�(Z6��1���wC�Y
�0�P"O�`gT5Sr̤ґ��2"O������,S�\ ���&Bi���"O>�P'@Z���S����\2�"W"O�12p�P�wm��@b'<1B���"O�I��Y" �bE0�aU ���g"O$=��+;T���1ǀ��qx�;!"O��׏�E�ތBt�לP\���"O�0�#<�� )�Jó4d���"Otxi��&��m��R�dz���"O�qBB���j쬹���{Ƹ���"O�(� ��(2fyyfl�A�(�k#"O�X)#�%5�0;�l<Q�$c�"O*0�3�^�w��P�(]�upq"O$�u���4
���6!�l��U�"O|�"�k�!�aa `L�>��Pr"O~�� ,�$s���+��E�O�M��"Ob�J��C= �3�A��9^H�`"Ob�8F((�e�� *`�Bq"O�$�(C9�|��m�!� )�"O��9t� _��sGB�uk��iT"O�!"BeT=��)x��W�cH^��v"OPy�`]��6Лbm�*09b�X�"O�ѳOB�/�x�M��:���"O�;��K?Dm�*��E�<>TX�"Ol ��#�.= ���q)6
:��"O��u�C���8	�)ں{�"OF�Iw�%��$�Ȅ�EĶm��"Ox�h��q�Ћ��4#�V�Ag"O�U;�lͨ]�:]1"�@�,��"OV����:�q�4��D�d���"O�t�Qb��jp�eOT3�&ж"O�s���?B�9W߃mb�9��"O(
&�=�d�Si�8|@,:�"Ot$RD��j�	�� r�2!K�"O$l1���%	c��F��H�����*OuZ,KN�t���*N1n�`[
�'�<�#p�#�n�Y�NQ3S>��'u�t�B*��u�H���DX�\5�'�\;gT�gt� ��P��'\�(7N�1	�����Q�L9"ӓQrZ�c��K(���X�bq��6XN8�1�JR6X�!�� ��N����71N�Yb��f��'0J�q2KW>d�
dF�d₰A�x5���C�@�%�J��y��4|$ڴr�e��1Ì����Z!o�Q��ky�'��h6�b?OZ���+ko*@�Ն^�s��|H'O��81�֏�0��Q^�N�5���V�kz�� H������$����a�� 7�d�GZp0ay2� Eb��X���54��d��M�|Z0MR�t,����i+!�� ��A� D�>�̥p�J�e���>A'@�O��Y� �9*Q?SB�-K�9��S�M�n��j<D��"�����C-f����q�O($'d��A�OZ8���er1�1O�	h���-��e[�[�#+�8#O�X	�6`�
̢Ǩ�s�hr ����AS��A.�� �@���AK?f&@J�̞S��቗
]��Q�Sa�(�R@�OHh3!��5'G��"�^"LD(�"O�}�6��P��u@FgՈ
���Q���,����)���H�3�ȟܜ�C���E0������L|#""O�U�w̄�8y���q'�<�^鉖�ܧz�Hʓ=���e�[e�g�fEh���@�T!<11�Jt��gAd�5M_e�h�� ϒh�n�h�+_�U��M V����'�";��z�@'?ax��Q�5��m{J�0k�քsD+OH�ٖ�*SŊA3��<�E��+������+NF���&
S?Q7����Te������S�z�%n]����LG��d�'H1SH�`)̈́ᓮf�*���hܴF��D��@G6&>z�z&�O�=Ju�Z<�-ɱ�?#<��F�d�����	y���`F-j�O��@�m���J6'F�]n 0>|)�࣐<<xj�XA�>@�j�(]�ݞ�#�����~"�1�h���3)�K�BN(�ēgPr)8��P�����.�q�E���S�]�И:�'s|���� �FC�	���ȡ���h���׊p�,�S`A�=�� ȗ�vw`��-2=�Z���'�F��KO8(�8��L��S*0�x�'!�&�ZH��I�sk�>�b�b��g����9�訊S�G+`@�A��;��d���6��J�G�$DDj5�㉨l1,�SkĞK��U�)Q�QsrL�f<�%1��d�6��f��7"�x�o�lC��Wgh����`�O���O��?4���m^�.ef�
̬�����q�G�B�*�t�j4�+>e`MIq"O�I�AbVM�zx)����/PD���.\�&fA���`M���2E�9O�q��h��¼>� �
��)���*��7D$$�(�cD�)�����-��e�}�ȉ� ]���f�ÿ3�d��/�X�'F���jV%)k>d�B$W!'����Y�����Ŋ^�n��������QzD���	��ty��^��1��x��e͓�0�'�� ���%5�e&�0�/�Z�I����"aL)��`b���{��}�y��8 A�ϻ##j����V����J"����=y�@�����v/LX�oZ(R�*�@���((#=I�h�:� ��4��[(�1�N�1~�z�CЂ| >C䉬~�Ęb҄J�&�V���Ҙ]�7��PD�xyU��+��)��1���.��X�JϚ}�y�:D�LZG��C�&PKC� m�䌢�Ĺ>�ga�ddA�t'4<O.�����;��2��\��}
E�'�����j��]�-��l�$��		���"��Arh<A�+�Ҷ�Ó&A��H9㥡�f�'g>=�Uk
l�����j����@֟$�U�[kbx��\���)��"OxR���DI@�zc�ι �8�!0�i�l 1h�
Tid�m�(OzX�	]R��5&,W�M%�ɱ�H 02yjpϙ��yr�@�Ha����ܴ���2�ID�QRX�d�?�Q����)B�D�	����(�R/�U�T���&���Cd�W-��>ID�]��X���8���G� 88�<�M3R炖~�(rUD!|O�4e	"�a��	��j#�=R����'��ѵ��_jn���/qƁ`�F����S�I_nC�	 M���҇H]�,�t�Q��\�v�b�p'ꜰ c��Ӌ?���y�,G�d�`�v Q"�.B�,is��wB��}����6�̖.����g_�z �ѧO"D��O��ӂ`(u.�T���Ռ`��mK�"O%a�n]�Lq��DI]�HE���iNֵ���+j5� ��	�#���Dƃ�GR�t�&$Y����d�l؊8��`��?ɣP2ΨH���:6>�J��[x�<q��йd��e�S�7R���wb
u�x�FX���C!�,!��l�4*�d �"T�T�LJv"O� ��C
�����"�:�*���~:�Y�{��9O��jS�H���at��t�f�"Ol4cP(O3S�
2B��:�DPd"Ob��C&�oj��Kf��Q����'�(����_y
� �!��e��M���1I��z��)��"O��Ō�xT��A�E�lt��"���68�~H@�5�'%%V��@�+~��`E�QiZ���B���� o߶Rq����E	��PT�ۼ���'ra��𙟨*�#���Z�aӑ@�\��8D�0X�Ƥ**�Z,�h��h����W8pd�b�����|�dR�Un�(��^�)L}� ���0=�!OƋ�&\;P���D��+C��(����;}�):��4D�|xB��&R���q.�W�N�c�,3�	�U�Z�l%6Q?mXp�Jt�:G-��+�l�"3D���`/B
%P���q���� ��Y��
�>����c����ûX2\ �.�B���@C�iz!�ă"KN�A� >9����/[�Br88�dd^A ��S�:a�pfC �� bK�>+��!���!v`�զ�G����p�� v�M2?����i!�؁6��1�v��/�9#�M� qO��vHG	�"���Z����C�-��6,�E�<�V 5����N_!-�`�3Þ�m'���{r�5�g}����@$�7��U{X�+��y҄ a`�qy�LF�0���Q�eN"�y�DH�L��xر�ӓX�8�G΄�y�H�T��X���/_�\�S#��-�y��	�ʞ}B"�I�`}X2���y2	��SJ���l_aJH{�F��yrgR7$PZ�)_��"ݺ�/̓�y,S�gǘ���� �Hn
���E��y��B(a9���c�O�x0x�Г�y�`�Q�e�r��a0���"�)�yBm�Hc$\Õr	H
�-�y��
��X$F�)RV\�E`�u�����o�2\����h�:%(a��H�b�ȓ�a�fC]�"�n�"�<G����ȓE�t��TÇ9��ܪ7�T�]�ą�$
a�$i°~�j����1!�p��.�(q�Tk�&0Y3��+���Sd�!��*�� U�����E�o!�1��!��)���0m��ؔ��7���ȓC[@��A�{�����kԶ1a(!��y�(NO&P�#c̛1I�x��S\N!�%B��1%*����K2X���ȓS;���e��G�H3��/ 1��ȓ)���E�X�lS�4�p��y����ȓ�Z�!L[�OD�$"T�J�LC��ȓPֺ��q��U%�A�熋5$���ȓJU��ś�k���'��6e����ȓ_��	�� UD�P���@̑�ȓf���F�IW32%x�M� �\��m�ۅ'�,�[��#%��	��6�^a���	��7ኀS�>m�ȓ�@A欆a4�`����nE�l��|�pCS�Z1�R�����M�v���*8��e�xe�Ae��p�ل�"���p �XUabL���%J����`dapf�YR�ӧ
�=2��ȓp0�e�5���s�E��.D!��ȓ7z�dRv]�(q ���C�9��L��t��-���Pc���Nt���l�I&��)
H�ĭ١v�(�ȓׂ����ܹ ıkGk�]e�̅�4o �1a�
K[�����w�Յ�ѢȨ@�K�p�ճ����|	�ȓ	��S���r\ݳ���m�4���[R@ pH�"I�@+Pl��iFy�ȓB���Å�3�@����C����S�? r��SjA!1M8ɪ��2&�x�K "OԤ��E#�z���7=�F"OfX��i	�h�Бc�͒*;�Xb"O-Z5ə��fm���?�%Ђ"Oz}�v�2a� |���N�)���d"O:�gF�jfUY��-}$,1&"O�3N�T�m�L~(��"O\�bgLU�zT�t�-�y@c6"O
�3ag�)@l�FM�#`vh�"OrcQ � w;��k0�V6b��a5"O�ѡW�۪G�D���e	>�P��۞}������)Q�����?��x �c�G��;�W 8�!�D�[�I#BMZ0�A�C��W�!�D��6��i�A#eBԝ)�W
73!��ۆ(����d"S	1Z��)؝!�dJM7���th�('("삱�_+�!�$W1v�D	k��'{��� ��g�!��)�}�0�>�ٱ&�/{!���$/�D�!j�O2A�Щ+w!��W�� @�F�
������Y!���w��m�&a��F�l�o	�tI!������)@NM�&^<4 T,�/*!��|ʠԲQ-N���h�
B�I��L�{`��5i����G�K?tB�ɿ~4:�!w�)u�(�ŪQ{<B�G�л䘡s# <�##ޔ6�8B�	�8<
'ެi�D���B�ɭiԌ���A�_ ���"Άp��c��E{�����.
`�`Ga��f��bs)X��]E�'9�N�&��'��Y$I �2�OX	/�b��46��%���&x{�C �Ǽ{��P�Gײd�i��g>�	�2�a����03X�&%��E7慰@��9k�'6䁸P����p|B7��ij�͡B��ly&�g�xR�ԝ��H�y���Dv�!î�/:M@nL���L;�>��~���ȗ0G|�Wj�_�<!7��u��Y���Uf�噕�\]�<ɓ���)F��pr�
�yT��i��a�<�U�Ռ5��H�0MN�`���+HLe�<��"Q�	�pd`
Ī 	��p�U_�<q@.�!A8��SbR�a�2��c�FA�<�SO�y����iT��J��7b�@�<�G-E/l��Dm�@�|�pC�e�<I�>~���E�l�L�"e�Y�<yVE	8�RŒ�A� ��xu��T�<!�R6C|4 ��5j��1p��P�<Y�HD�-G(�A�̗	{��DR�<)����I�&�h#(G�7��+���x�<�� ����JF@@
+KF��C.Vs�<����u��Tg���2�l���ǔq�<����4K��̨��"cԁ��'�o�<Q���V>D����J�.�\����i�<q��?!f=+gF7S�@=��/�!�D�N� Q� �S����M�"�!�䚶%����B�ŵ���O �!p!�$�zv��䎹_0p�t�Ļ �!���9}P�!U�D�C8�i�bĦ�!��z����j-j���۰X!��d��̪�oB
��AE��,*R!�
5(�0bBn#��iG$Ý,�!�E<s���B�%@�2�jzG��9�!�ru(�I�d$J��{�Aڊ=�!�$��ki���%v7���f��d�!��y)d���@/���?�j�'�(���σ o}��G:�*(��� ,��ɇ�v�� (�?5��Q("O��q
��of�qp�ƀ�\�3�"O��bk�
�T�C�ł�'4�[7"O�򄮀�n�V��c��V�.���"O�$���$`L(�׈-7ϰtkc"O����rtA��'W�j$2=ѓ"Oq�7MU,0:NdG�7;4ޤ�"O�lȕ%�.M��$$aS�/4�9�"Ob�ʣ���`��|9Q@�E#���w"O�d!�c֞���a�m��""O�i�v/�e��t2o؋�t�E"O*�R�ڇs�����N	Q���r�"O ��Ǆ�:D?��y���0u� �	5"O	�wC �#7,T
T��Mӕ"O^��X�q�T#P�ϡ�Ӈ"Ox�0��I3/�T(ۇ����=��"O"<9&��4l��E�3,B;�dt��"O�§̒C�Ȍ!��O�{���A"O�8����M�Y�E�	���$"O�4���kv�7"�p���@3"O�=�CN�Xq°`
l<��7"O��ar% �e�$�R�̓%l-�7"O�p��ȃN@I���A�P:P�"O�-�DFE6#�+��Ö45�"O>UP��Ԛs���-S�]�8�"O�ԊRV&���ғa�Db�Ic"OD�:���=c��0:2,�a�"O�Y��H�f�N�r@ɕ
ɸ���"OP� �q�P���YT�AS�"O�E��	�[YX8s����eh���"O�'\�W���a��+��`"OR�*E��Zb�E�ƦB����c"O�����,~��3�5�h�P"OX�O��DN	����
/r$���"O��caf�5s�H�ݻC<�xe"O��I�ќ4F x`*�Q2�5hP"O��²NJ9U���Eʈ=b��S"O���Pꚵ%�.���T*��)c"OXѐ/��7��H�S��4uᬈ�3"O�d�c�)�h8�V�߹H��Y&"O�=�ë��>D���?���[�"O�H�G0|�~A�Q������"O��H!.�-ĕїdTE�P|iG"O���F�4.}V��cѻ`���a"O��R§] S������$�(���"OIk%� ���{�B�t�}1�"O��rW'P��>}�!�8*Y~8"�"O֙�#fČe*��U��<m�,�U"ODl�4�Ԡ@���j'OB�T��9"O.9S�c܌o�\m;�a�`Y �"OzzU�� |���Ë_��j��"O����	0d2����!��	�h��"O�A#����G� `����.n(��:v"O�`ʰ���b�b��F*"~!�"O��)��Ήe����Ċ�s%��"O�؋C��4��S���]e4I)�"O:�F�x0(бe�xpq"Ov���ʘ&�ΰ1�ͺ)K&Md"O��t ��\�&9�
��0�9�"O��Y���|R��
 	X4�q"O,�i BM�,Z2�u�����X [�!�d
� ����'�9�A�p�!��»��(�W��J|�ԁG�.�!�ּM�������N�@b�a	6@�!�� $t���B��0Ph�
{�,�""O�i*`"�X���0(�k�<0"O~�I�3��q�&��o̜e�"O�
��ɯ���T�Yj���"O��J�W!r!
���㕄 ��Xe"Oƈ�����J��6�Q�%��4��"O2�"#D�YԒ�臢��Ct�D�Q"O�]�%�/��1�.��.���"OP����g�����I2 QH��"O�ݑ3AJu�~5�כ�r���"O�=闏H�Q�fD��A�*v���"OT)85Ѓ@u t� �=JsP�a4"O�Q�����Fp0��vO-$4["O2����
[$lS��:^�ص+""Onh��k�iK��`��/q�r
#"O���׃ v�NUJPΓ�ֲ�QT"O�T;PCA���MD��Ns�"O�M�Ć�5FG�y�c��UQ�"O��X�ɐe��`B��$o����"O�)����yV�`!�h^���\R�"O���q�Z�6�nEcr��Gġ��"Op���?!إ�v�D�>���pd"O�a[$�� *��q8W�	� �*-�"OJu f�I�m��h��r����"O�1��养Z��	Q�NI�z ��"O����\�A"R=�b� �br����"O�E�#L�'>T��K_�8u���"OD5���Y R�<sE��lW���"O.��a��ָQ���/q:*��"O����"	/ �� Y�i�AC��"O"�w�ش:l�2 ��?����a"O��0�\�}"C�D���k�"O@�����z�A�6��t����"OT4u�B�
���qO!	�~%�'*O��	���/� �ж�կB@���
�'�愣7�aj��J�"���ܴ��'0( ��^L����-
��<9C	�'Ő�%U�b���0�u����'�\�hoT.ΐ��;x�3�'J�DM�*98M���		%Ȅ��'|SUJ�	-�xӒII�6��\�	�'�0=���;D����G(G&d�[�'�EP�F�>|�TŲ7��-a��h�'�h$i���u-(�P@�['NO��(�'Ę�J@B)씪����Rw\�Y	�'�d@�4a��vߴ@�gL�$<7|��	�'��M����큃E�>�ܹ	�'ת�:0�I{s�8�eWir����'荃w�Q�6'XM�#��c���#�'��ѳլK3�J�aV�	
Vi\��'�|�(��<c��iC��|�9
�'Zm�GfA^:pi���-4R0H	�'�J=)	&�Z5I�eF�[���'ϮX�A��3kL8`҅�0΅�	�'%BI�4N�*���fC�;S<�	�'�$��@QU�vI(f��<_�L�X	�'k ��1R�Jdg앻.P�,��'P�,)�3L��I6�ّV�lX�'H��&��'Z@4�6K����ʓ)���{	т>����c�w��Y��d�3[,��p+HZq�Q-�y�!�.pY����2oE.���+�+�!�đ�fn���ԂɬE��9��N2W�!���.W�F����e.��6NX�Gx!�� Vը�L�'`��rt�Q�-�܉h"OT�iw&ř�a`agl�M�F"O�Ī�.Ԑh^� %��/pa��f"O��h��^�;�X���Q+%J�4��"OX`�5B2%1�8��j̚e��};d"O0���L
� ���h�_���!��
���Az��V/Y��-���J,.�!���r���_7�j�����3|!��&=I8;F���X �1�	g�!򄞔,��p�p
�X�����bL<>�!��.aTr��#��0m�D��@G#�!�T��*�p�����1�gL!�!�$O:p�x�$�$Gf�͓��h�!�D�QFJ�5� ���!�ǝoi!����ٙխ�~i���`[��!�$ӄ<)�4���^fL��ƙ�(�!�KpR����̎%o��������!�D'A��D���hP� P6,�!��K�Q'\����"RҤa`�W6�!򄀁F�
�(�+��Y:��S�͗r.!�d��s�UZG���a3�A�2,!����H��.o#��sg�#=�!�	�O��aH�@�30�M:�H�/�!��1����F�(	>�&fÒ�!���6�j���n�g��r�EO�/�!��>|�� \1z������U�4!�D�"g�	�$$<�d()��ůc�!�V ^L�s��?/j���`�`�!�D��6���bs�Q�,L]��*�	B!�dVi�y���՞
?����ީ"_!�D�x�z ���j.��;���m�!�D�)�Dbum��")���X)!�s\ x���7?2�R�1J!�d9wq�1(�=<��³�K�M	!���I��V�LT���+�"H�t�!�$�`?,�� k��N�.��D�*�!�D�H��L�w�A:�R����:�!�A#�N�:!ʓ�D��h�)	C+!��L�d#�!�p Y�f�B�S5霮,�!�%1j��@�63����G�����9Sbx�'��O�q��D�]]4m��o*F�踠f���ĭ:��Ͷ��˟,1�O�s�'�"�ic!��r#�0j�-���it��pyj�D�8��d{����س[J�H��ܮ2������<�rd�I˟�:+O��:�\?����;k�V�QQKڷ:�.��A)�68�����'�ab/C'EN cf��<����j���d�<�㬋�KA���|�'?b���i��:�mո�
1�f�*���[�'@�����+p�OBxQ�Ιb�m�>e�Blߔ*��|s2 �X��������(��N��p>iN�&1Υ1��ޝtc�A�Fb�2ѫ��3�>l�Ԍhi摭;�O<��!iI�9�d�en��`�1��S��P��Iߟ Cٴ�?�-O���;��f� D2��,)C�TrЭ��n7Q��DyRB�<yc��m�A�E �b�F-��g��K�6�1�Đ8K�n��<�Q �B��\��Ȅ�w-�+J���#�S0#A��4j��g��	��\��I؁��S�S�ȋ���]��1!����C�H��CS��c�~�� J�(& P�;���+K�`�]�:�t-K!g٢���r���O���C�e��`��@!]����a��%�|�l�ڟ8�'�2Y�<D���>����E2,�H��X,�hO��F���iu0��t��Y��]�P�@8i~�� T'��qu����O܉oZbP�hr�E��ȗ'�����f�����J�"r2h�C�)Dt�J�K���y2�':r�Q���Dc?%Bcg�����Z/k�� 8wC�r\d��V���k�dM���F�X�b���@P�?��O�U{��	W�t ��m�%
� h�}bAI��?A��-i���'ىO=z�$�U��<�B�*�,`�ӣ$��"|r�O()2��,W�"D��暁0�ɑ�'�6͝ئ�'�~I�!������Z�DA�s�>A��H���@v?�+O�ID1k��b�(�c�"����F�3<oԭ`�#B9D��А��	�<���fh�(��lΙ"�xP�?� �L;1JU�0mZA#N��I��±a@�!���� 

��=:7��0�F���m���M���˗HM�B	�1bf����?���t��v�'ʎG��O�-ũE#,W�0�V��c81)t����T�	R���OQR���;;e6��s�>(g(�"*O�aϓ%�f�źi+�'�뾰��֦�B�h��w^`} �-���� W��x31��>�N�?-�()����<I�4~8��b�Ыz�܉�7fSU5�7-6d0��S	�+(����V�L���+F����!uL��7f>4�fI
,Ҭ��s��k���pAAn�#?q��HdO�ܒ3��y����t�Y����O��D]��T�	q≽-�L�+� B((ܭ\W~��f�/�O���'��cGh �:����� �6L�f1�b��O �Oj�(��Or�O7=�lxQ�  ��   �  b  	  i   r-  �:  "H  @T  �`  �k  5r  �|  �  _�  ��  �  C�  ��  ��  z�  Ҹ  $�  q�  ��  ��  :�  {�  ��  �  ��  ��  ��   ] 7   �' ^/ �5 �; 7B �B  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf�x��)��2���T�)��A�bV);�C�	69�2!�����@���#7��#=�ǓY�&�jE�B2w`U`I(P�8��ȓ���Ǐ�FH��{Ѫ!]Ǫp��<�L4Y�
Ɣv]��ٽ2|��2�	�	E��['�6\c��Q\x�� �bK:��<���	�W�T�!ҮE�q��L� �2���O,�=E��I�/6�����
nO��HDcV�y�I:?<��Sg�j+t�@$j��yKJi�1� �
�3�T��3F��y2+C�dϦPyI��'��Hc����y��'��D��ŗ|��e�h4tTyS��D8�mH`̃uF� v>P���FH��P���Zp释�4�zM܁\R�����hO�>]�5mR1NX�Q	%5�����>D��
����,ĉƯ��^���著4F{�����d�+��J~�P�SBE�,�a}��>��(�\�Q�Ο;2�P	��Qu~�
)�Ov�G�O�W*ʍrB��K�rR"O�Csc��+�ʌ8 �k 0"O��Z%�,��d��M�*j���"O�M�"O�d�1qvj��kj�t1�"O�t�F�-<Ḓ����m� �"O� 451fn�!�N�r�N`6ޡ��"O*}�JI$jy�H0@ȁ�"OČ�� * Pq���(��k "O��ӣ��2ۖ��c˘���"O^M�c�"[�ΰ�O�"1�����O����@"c2�� �.���*�H��d!�$%8miW��lI�Q��9�!����k[x5Є#�%R,��;�.��O̢<�J<�$���"-�GO��x���t�j�<��B��ؚ�L!/�yBP�p}"�xb Y���i�$OD5�D�A�1g��Q�*ϘO�az��i�	&��7b]&_B���
88�0^��hO?�*�\-��&��<P.�p)�eqON˓��O.�S"l(���i�Z�d���ЛP���+��y���/^hyA���5��SF#����b�>a����I�E��Oc��r授e���e,��gG��s�'�Vu��K��gMVI�,iC��)�'!0��ȂSd��O����<�����ڏBLM(0�I�φф��M�UKI�$٪�1��=�D�*�eP~�<�F�FT$�Ibc�(A��!�AvX��Dybi�:��p���ܦi��GZ8]�F$���>�1�H�+��i�'@ًt0~��m�	r���Oo��,��2�^�>�p����ؕ�yaR3 �$Hf�ͱ1.Jp:�g��y�
)LT|QЅA�=X��H��y�M,ls�TA�	�^p�_�8�@B�	�lf!���ět�t����tpB�	�)��s.�> �hx�5m�*; B�ɺa�+�*�+'����+�8�"?t��F!޴�B ���t�{V@B䉄<`���\w�A�aͅ]u�C䉺�� �UE�9~�@�0�~{�B��Y���`e�Uw���"��NB��S?��]�N���Y)L�S�/�;G��؄ȓ9ŔmZpc�o��af� ����ȓGb�ñ��3���
�oIux��ȓd�����fؖ?"�ѕAD�J?�=��'b$}C�BO~�h&#}�����f��a��b�`������ȓ8�B�h�oi�2��
�&����@5�I�iˁI��Q�hS-tY�ȓ?0���K�,�\ q�KP�=>��G"D�&M0Jk�p�Vd�!mG����Uy����Ϛ% �)4aK�b�`��ȓAe���ԥ
?�����ǃ"o�D�ȓq��� 
�E����`�:V��ȓ	�2���nmf�9�S�K`�����1�C��6Y�.��閥%~���s�($����
� A���i^�І�M␨�`�=����K"'�ZІȓ)�&�Z�e�>u���@�'�`�����Wĕ�&��: ��⇻i�� ��8�xɀЁe�fՒ�k!Y0�1�ȓz�͒�A�%R@�ybS��\�l,��w0�9����iH�m��!�:O�9�ȓSN"�C7-�	S�$ܫ�ʁ3k�
0�ȓPO�c��\�c����Ӧ�\�Z��%��b���k�"�!)��I#���3~|YTaàT���P��X�����|9rF�L�o�4Y*����ņȓ�0���\d4��TD�@2�Є�B|I���o���Aʇd���ȓ2�x���F
,�젩�l��D)�����l9�$��c�ɈCd)H֜��S�? �%�j��7G��)	��S���S "O���ŧӵ[��0H�Ʋ���X "O�劆�>2��XA� 2zF��5"O8�˰!�wN� ��e̢�ј�"O<��Q.�+9,)���|.��F�'��'>�'2�'L2�'vB�'��!��ȼCO�[��+;h�QRd�'�B�'F��'ar�')��' �r��xh@'͹U�p�S�PJd�P�$�O&�D�O&���OJ��O,��Op�d�O:L�5I�j�������y@�fg�O�D�O����O����O����O���O��YƥԙlI@�z���b4L�RT��O>���O
��O����OX���O����O���%�t᦭��� X�0bG�Oh�$�O��O��O��D�O���O��2t�N�q
�쒢��n��%2�&�O����O�$�Oj���O��d�O�D�Oz��Z#Ŋ�c�d�Y��ܻ-�ON��O����O�d�O"�D�O����O4���^h�p���&>�C+ӹ�?���?	���?9���?i���?���?�R3d��MYg��3Xg��{� ���?���?Y��?a��?���?)���?��@�4f[�d�9Y��Q��Ԅ�?����?I���?!��?���?���?���xt�I����vZՑנ�?y���?���?	��?���?���?	��R�NL�M�V���ABa��L#�?��?����?����?Y�������?�nU�Q �s�"o��!z�j�<K�B̏�7�bE��Z���'��'�6��4�,�q��A�V���K�ɘ'��6m�O��S��9O ��_);�����V�mFH2���*0|��͊n0����'\�z�j���'cD7��uׁ�[��ɱ<e�q3�\�����5�ˌo�x�a�4�����Ȕ'��fT�Ӟ�XU��*İM\�⠇čK�l)�p��[*6c���3��Mϻ`�&�8�!ф-rJm����
���?q"��{�BgS�v⬑�O�b�i����I$!ߤ�+n��{����I�HP�'���e�^�8���1}24O�!�X�?��]p����������#b̓��7�D�
1���`���~n� �ȧJ��d��������������O
��Hc< �I�?����4.�/)���А�rmX��'��Ʀ}�P�
v�(��|��mH؟,�r�w�v�AZ��j�M��O��)�]���I�}��8�%�&�s�<�'Ȃ�b���t*��4T�q:�����'�07-�OX�IU�I�'@���ӫ[��y��g�x��aY��:�ę'
/�����sݱ�'7�؞�u��bW�I�0)��9F�a� ʝDRH�*�>���'�$�@�'R��'�"�O���K�:猀��Cמ)���ba��	��EN��ňNşh�	�����8BY�'�~!��$׬WǾ��$�$x>j�JE˼>9c�i�l6͆�i&���5l͸͟�������R�!��DҌ7��@!F���Z�4�����6hF�Em�a��C�>O��� ��	�?�jҥE����!�	��s�V\���"��?���?����?q+O
ʢ��?/���'��(�́5C0A�Q�G�r��Mަ-��A���6 ����$mڎ<,v�"4��uϼ�+ӈ�0=���Ү�.|@0��*?��N�D�h��mޤ���T��݉v�nIQ��.WT��8�d�^��%j�ԟ��	͟���?8V#h�sޙK�9fߪ0�c�EtG�1�����	П��6�Q6[�J���4Q�4�?�2��<a!h
��iq	M #��	���
����x�8D�E�Mϧ4��`	M[~��T 02�K���C�h�5jQ>+׈�r F�����`�f~/�O��P#�������?���u�8�j	�%�4p�D�ё�>�+��?�*O\t���
8Ek����O<����Z�*yCAH�rp �$7.9�ɘ��$A��� �np��	*��x�r9���Вi&xơ��	�.x0̋�(i����d}	�䀢>��"|����#��L`tH{ԡˮDb�Y����1*k���T�'2&X�r��)�����'b�Q�DQ`��&<(0 �43�Ѐ��mʐ5\�I��L�I��M�)*t�'���(��Z�x�8K-R+2��(&��b��7- S�+��]�&�(Mq&I��D�#_���Η=ZR}"��N�W`�2v��Ou��)~M�q�����	ǟ�S�I
x�O�����!�[f>�CsF���֑�c�J/b,�yV�'d��'���'f�I5�M�;��}bV^k?����8=�r���?���
]?9@�L���(|8��]w�ҠٍU�:���̌���*@�
V�󄓽3�<�'�zA�O���	7(��'��[��P�e�� ވ�8�ΙR6�' ��'��I$Y4Dz!��d��Ο��W� �f��F��~�2����V�.?#P��޴ ܛ���~�C�$�:����ؚ��$xǮ��~�THΓ�?Q��]9pX����J���ú��f�꟨���O��4�A�		��B 腖Q
�Љy2�\Q�:�.���;&f!�$��z���!���?�'(�M��و��?�b�i�� ��4�6��B���RrCN%$"�y�@c�]�x�*��Q����g�ZA�`��??����d�<֝�.��ыV�рh56|�v�'�6l;��SK�C⟸3r�g��|�D/� G\�0{��]}�d����/M�ڱ�'ˠec����R���'����yʟbYZ���=����%�P:��s}Ho�Im�J����g&,i&�?����ϒj��I�!ϢP�8:��P�n:V͡��ۥ��D��1x�y���T?�ѦO)�	���8��5MO@��Mc p����T��d��ڟl��џ��	ay��^�	��#�'���bZ�.���b��Hdq�!�'!7M�OV�� �����O�o��MG,�CA��C�t��ò)O�E���������nZ]?� K�L�]�l�vᥟ�	�=� D���IQ�OO�)҂�3{F�+�b��'���O����Op���������Rq�tR�
=n��C@��]a����O��dO���y`6����J����p
牤ddlh�G084󵠐�T� AZ���\��ȃ�0�nz>i0��08��K��� ��	S���փ
 >�1Z�OC ?b���۷J �?z��G�R���'���'���K��F�Y2�}���9���S�'}bR��B���	ɟ����?�-�h�SႄZ����nW���	��I՟��I�?ؔ�I�E#P])70��M��F=�t�9AC�]�"��Bo��h!B5!!n}�\P�O����y��d�$�.V�1:��7G���9r��4���I$>�t
�
�ȟ��i>�����Ĕ'�ڐ*�K�4s�2�a����M
�kto��?��O�pm����q�-?!RP���":V&���1�X��6�ȏa�����2O@���7˂+`y0��ʟ�S`"
���iF�H�'����-̻
~<��E
$d1�y(�`�r��/��'���'k�D�Ch$�Em��� jZ�Q�v���g�#�����$04,�I�D�I�?c�d�����u��UH�-���1��X�2ԩ�?Y�* ���~L2��;z��,�u�4O�yt&9!f�l��،��l8�5O��"�i��ybȎt��Lٟ��ԏɝx��	�:C�E�/ƴuZZ�C'Q��IƟ0�����'(��`d�O�c���'�bɂ�p�Ұ�7HK3C� ��Flх.�R��3����t}R�x�Fam�H����j޾]�A Ert6��!'4~P��:Q��|�O\9���%bZ��S�4�`��D>����5];�,��?P%�a�F*�?q��?�S�0�<A�L~��?9��eibxIwH|��53�׷HM��:�i'�͓�?��e0���'�f��O�N��R������x+�Y(8I�)q�ŶP`δnn�V��m@�4�&+��VJoݡap��|r�u�4���hX05 � >����O���I<H2x�����(��ğ0�#�p񪅨��lYp.��?������Oy�f�2?^�9�'<��'Y��ybm�: �1��6UB}sD"D�]הꓝ?���!ڄ�h�XX7�?�
>��{'gX){<X�R*�:m]���[6Z��ɖ�*��R8OTԒK����#�e��Ĕ�0��}��m��*"���&�Z���?���?�����@5HLx�5�O0Q� Ue������F5_n<(d��OH�l���<AP�3?)V��Iش�F��2���n<n�4���A>q^�[u-M>x��;�O�(�J4�u�H7fJ�'*��E�>��BCFۆi����n-L4�����'qb�'���Ok��#7���w�=�ȃ�$�ՙ�#-�x�b�O
��A61�1OAoß��	q���蜲������KAH�<<i@X@3�O69Xd'��O� �!��D�DΝ�e��!q������9z�r(Ku&@�OW��	�+�L�C��[��B�\������d[���=$�xQǌ�;2�	��.��D�	Sy2+D�y��y�'H��'��d�i�2�SѪʷS;R�����$C�`�����0�O��$�O�|#!�OT��SDܥ��cZ-Lς�����<d�%(�*2�M��eؖ��6b�P}��3z�u�h���'�4�K�g�eZpus��3�\5҄��O�my�՟��d�O�	�Op�ĳ<Y%m�Q�:�w�%f_�I�ҜP��Q�<��i��D�����n}��'�h�aD�2�H�+�$��T�у��'F��c�I�F���O(�!�U)�u�4+Ep��k��1��K�{.� q�$���0�ɼ�?1�
�W�FQ)���?	��j�/,����~7�Q�C�?豲�jB�m՞��	L�D�O0�����PT2���D���,3F	�v)L+2�H9T%^�aUvM��蟔"#ʲ�X��$�oO���E� I��+��2q֧j����U����k���yF+`�rϓ^���'?�䝼	Qx�g�:�*g�ݩT���A��&D�rq��	5;U~���
̟$���l8b�N��	��i�,U���AKƟ�J!h:?��V�,A�4Q��k��~�D�6{-�!�`J�G��$�dW&{�@H���<QTV"	QP�b��Ďp��%�OvhH	�>P���!�*���ᐫ{�F��Ѝ.TH�$�O��䇆S����4�,�	�O ���OQ;B��
E8{������a���O^l���<m�B�'T��q�L��V23��i���0eZ�=�*RDɲN��AhC��:�2��2�MK�iJ!5؄4c4a�O~�,L�B3�L�;	V2�kP��.4�Y��h�<%��ȅ(��	��?	𪌡����4�A�u#&e����!����.	������Of���c��D�O"����?M�&���},�lj�Æ07�������dæ	jٴ2}0��Q�B�+W�-*7�ֻ+��}j���5FE��(�܀5��(�`�݌W���Γp��k�M�O��!W�>��'�Na�b�[ ��8E���|xwdSL�Bő%�'MR�'Zb�'9�	�"��]ra��h��	

Jf��* \��������h�4�?�!��t~B��>�3�i�h7-ۄD)(�Hn� L>�h�×����`�� ���B����ɖ.���ל�OI"�.��V�Pl)��VNˌ�E�ݼ �N	�,eӠ$�	֟@���?] 5"Fj�s�q�l@�:[�������B�Z2$�� �����9p�O2�q���'���ț'��LI��7�J�����]l��0�N6�~"���6*c���t(E#,�H��� ��y��U�h�*�
�L~2�;�-ZO)ش�F�4Tc&}B&�O����f��d�	ޟ �ɓh��MB'�!�4tӲ%Q�n�����ĕ'4<�W%؋n�R�'����y"I�s�X���ɴ����N���]}��'��=�~BD
W��'8�D�u�7o ��G�<wD��#�A;zij0�ٴY� �������F2�&��{��i�Z00��i� i��M��J�^(�$	]H��Go�O`�4�Rm*rK��˓H�&�ѓnŽ;�d�8��X94���j��<�+O~���OJ,G=OL�$�<)���@y+�GA '�^H$i]�`�����^~ԝ`тJ�̓�?a��ع �X�۴G��S�? �=`� ݺx�T@���N�z3�'���DD;s���O��d�O�����O�L�'H]>�pP��i#H�KKR�wH�	��@?$�2I���?!�����|z�w��wQ�܀�:V�����W����'N�1�~��0v���OװM�g����P�-=p��p�S�*#NکA�O�7�I�'+�:�4OacK��;��.���O���]=/��u=E���BǦ��:�����O����O|˓s5H��Eʶ�?���?qAǂ�l�n�B�C�B�ɣ���+�?���T~R��>���?a��L?yq���d��x����!~w���i7Qg@�C��, �+��McPM$�D/A.�y��nր�)��`\8qQ2��hR����O���O������2�����D�O����hOT�+�D�4�*��eB�46�DC1
��$�O��R��m�I�Z\��ӼK�I�"[����	/$�E����$�v��H
���­u�U �@����ĉ�?�.��Yw���k��$2�58Bb�~ifA{&o]2b�N�2�
����'[�'�����xP��0�d[O.UهӧZ�Ή`�T��9�N�}�q�Iӟ���?�)� Ƙ�O���z���L��q�vc��
;��ӟd�ɶ���	J������?��AAO�����J6��2����}nZC[���$�<	1>Of��n�<i��'�����B�R��S�mޏa��DhDL�t�'��'���'��I �<ᒊGן<��
Ud�6�+�
����%x���ܴ�?��H`~�>���iD&7�H�N�93p"6U�\��b"��c���G뜯�5�����;�?e�٪_w��OK��*H.\@��9tJ��0Y�0ۧ��O����O��D�ZxB�%>�9�t,�6�3�XɰLg������>9b�'hr Q��yʟ�<l���Ir��q��Ú��9�f�� �}���>��	5!I<�I����	�ӊ.5 1���O�|��b�:���@� lPI� �"=�&M�Z �G ���I��?���q���OH�d�O�pQQn��[��->S���S�o�Ob���<Y��A�Jw�����?����3�L�6�Q�S�8L˂��(mu�'�8�l�f@sӺ��3�O\��@Z9��ĊSM�f��&P�I <�6O^(H���4kR�N �z0�Kv?�S�U�T��U4\x�M�L<0ECS_��q��K'�n��'��(���0=d��T!(�@u��P����ΏA3��jb]	�?����'��z�O6��'6MS4y�� �&�R�JP.�;���m�O���{��7���`�O8	��NA��u�F^9l6��,��`�%<v~��`h���~��R��y � � ��ȟ��I�?Y�p���d�AH��*o�n�6�:�b�[����/_���'"��OczY�͟^�mzޙ���|l
 ���D;%[ P�E���MC��i��u��'+6��P��r�t�; Vp1�eޢt
��!Y�J���ө B�=��'O�xh��ꟈ��`1}"��O���O��$�P�����on�$�Ą[�P����O����O��3Ì�i�MM��?���?��)$�l�4薆]N���P�?i�&�Q~ҁ�>i��i����~�Z���������u�ƍC2 �'9�y3��Jkd<�5�!��O��?�F�|	�A�W���GbJ�\����R��O����O�H�#b�rp������O����+�r���e�Qc�]a�A��
x� #f:�$�O`�Ć��!��z��Ӽ����1W6�	Җa��?�(�a.B$( �y9Pŉ9m�� �_>U�]w+���h���I�"��h8h}`p�ߠ"إ���H4K��'�8�DO%$a����O���O���ʹ4k�9a��:�V� #	C.i��K��<�p��&�����?������|��=�Xs��ݸK�	:��%�z��C\��pش#�2I�O?���	�ζ�>��)�S!���hIR� �v�Ip�̉JL��%[�P0�Yh�J�<��	�?�T!V�fc���Q�}:��)���+���hG+���?����?����?)-O�(y+r����՞D���R&� �J8��r ^�Z̦]��)Z�J�hh�Ɂ�M�q�i��@�0*Ex��3/�	k��A-^�r�JmqХ���ڛP�z��Xw4$�9�~��w���ڔfS4s����ī[����Kh��'���'����]=q��y�
"Y+��[���;2���j�����'��"�yʟXn�����f�{�`QC���+̕򚀑"C�W`D���FL��O�IN���T�ոi'���@-�0��"@�Ģb��YYf��M���y�	������D�5�u���?����?���T�I���3O��`i�%��?I���>��h��g�Of�D�O���i��S�NO+���*���%l�hO8?��Y�0����-��Ƿ�H�����3����kl\��oŰ1j�%�e�$���c�fڗL�3��܎�~��Iɸx��C����'l�-��'Nv�h��X�5��4�)�O������K�.���O��O��ı<���I/
�(�e#�0t����aŨB���l�B�ĂѦ�I�MP��I��t�����S�M�8y��L��� �9�&�(F��m� e��'й
Z�L��#^8�z��O$�(D�V�pa��HŃĮ_ \�6�'h���e�J�z@�O��O��)C��t˧M��CR��-f�Ь2���Rul�g���?I���n:����'d67=��(�FJ�*Z�D$��f*�d|e�Ҧ	A�4�D���%�����.���\8�Fim�:q���u�+`��sR�V�2p�'�a�A�����{u*TG~,�O�JYw�08��X��@i��]P��X'��wd����?Q��?�.Oؐ�*Q?X���O���c��рEeU>4�QzÈ�/1���3+@�I�����-�ߴe�$����E�)R�U�,�/0'�+1%ٚ ��I4bS2P���,V~��Ŷ|2����L)a�w ��Ā��-�fx3WG"8ł2e�'<r�'n�t 0(Y�0�O^R�'2OU�+p��3 �Z>�x�#��)��ќ]7�Ox�D������5��Ӽ��dΘHX��!��0*�iq�L�zp�P+ ����&�D��1ɜGL��'�u��,Y��Kb�:� LAw��u�]���	! v)xfI�
t,剑�?�6����Mc�'�2�'���g��g&�%���LA��R��P�cU����oB�xʹ����Qԟ$�	�?!�ߴ�?��v�~�� .�D�������i}:6\����4y8�&�t?9���!3�����?eʔ�M��t{��~�P��'��{!�+PЊ�	4��a�G�'���M�<	��'S(��o�&ls�Y�5��
�����'\�dު��b�'u��'\��'S�ɿd	�5��gK����%�]7 [2 �I�%��%� ��D��4�?ф�b~�>ђ�i	86�-(~>A@��B�U�$��$f�M��9�S�R3h�$�1�v<�̓awr��5!h�!���	NX哒̿�b/�&�s#g�"Ff|��u�!�v��ڴߘ���eӭ�O�i�^�<8'�	�X����O��d�O�0��F�զ�כ��'���c�'a���eՁ4e,U�r �zn��2ƙ��~R�\�K���R���t�8^.U��mC��yRƇ�
�	�gMAtH������N:JP�V(������������a�������?�v���a���j�p��$#EA�:|����?I.Of��2��"n��d�O4�$�:8����-a08"���&H��	�4��I���B¦a.�Mc�⺟����Q��)�$ux��e��;,��j�$�	�����d���#DNZ���O�B�9��;�v4��P���n7P�P��D�k}��0��N�?�T*� ^H1����?�'�?Q����d�T��H!c��*�h���#0d!�0+�ʦe�I͟�
ٴ�?٣͍F~�
�>ٱ�i��h$��i> @p�r*Z`&aӀ}�e	Q�i��lL���X�4p8Xw(����@�<Y��\�XmI*P�L��L�f�A�(���&�BP�ܴ)�R�'���O�dy#\>5zp`U��yp���!d!aa��3��e_ǟL��П����M�(O��mz��cw�фZW^$ȵd��}F.Y�E��L�I�\�:����RpCr�?��MX��sƍ6H��DZ����+lW�M�@	W�<�5��[���'�p��'�f�$|��ic���I�c&��I�;+�:� �P	K�a������ǟ��'����W$�<:��'��ƈ%n����%U���#�OֿqD������z}�"�:�n< ���	�d��x�6�C�T>6���Ѩe�¹�F��jm��S73|NIp�k�+o�~)�V>�!�O���;z �R£��PFyQ$K�r�ʈ����?	��)�L�"e��䧾?��-I��?�,�s\�r�	 #}��#醩�?���[�v��&�'q�xӬ�$�]��O�n\�Oo� �ʏp>֬s�ŇI���b��-�l��t�\��2I�=�Yk6��ϟ�� �E��.$L�����A�V`X[㯜B"�-Vl�:�����i������?����*$�͞I1�hC�` )Q2i@���C�,OƄY���L���OB���b'�z1˛���1�t��.B� m�riB!����O�����dͳs�:Yʟ�Z��F`I�b�v�v�9�ǎ*C��Uj�e���ǵ ����'���#�X���'Q�|���;'�  �2a�%̩)�ስ+Z����?a��?����G�y]�A2�k�O�8�W ��ϸ5��S'45�M�1b�O:lm����)?� P���44����Ɋ<h�a"�g�����L��4U�`�3�"�pv$Ԫ�y��L(q☭�H=�)A"�|:��w���Fė|���#P�º ���C,�#rE����OR�d�O��i@�g\����C�^h)pΆR�R��fW3 �&���Ot�dìNDpo:���i"�Ѵ�y2�_$>?��v��jt����K�%B��MP�'�\#W�G�o@��O�r��w���L�'�&���i���!�6&L6����� ��N����	�:b6d{(O� �ɬ=���m�#�?����?y��Ź\��r��}�v쒗i���?a���dX�꺣c�/�?���?��':3�v�h��� �M$F���ѵ��8�y�'��w�vF�O��[�'����ޔ��D �?	��*�KH�R#T<�`�(V���P�6���zf�<A]w�*e�Ͱ`Y#�OЎ�!'	?�b|�J4z4������3 ��*J���6�-:�V�ɑ5	��×�A"VW� C ��&�8�b�H�uF��7�֜^I
h��HM
)~џ`��ߡYuta ���3'���2ID�F� ��V�R^h���c����ى���pV�@$�?+^H�@蜘R�P�`��~��re��2�&9H��G˶`�"%	���<�)z�Mֽ3�&��S�_4l�3�!��y�L��Y.���hTq$A���Z�:1C��g�l�A���Y� ��U�%VQ�``�O,؁0;O*�d�6���O�B�'��L���mn���gָS��z�gN�'9�'���'w�V�`�b�I_��CS�#\(AQ�$%i���K�Lצ}��� ��b����"�$�OL��E��xk���r��ŻR"T (�����>y��?Y����D�*���O���S.JW&qғ�$e�*q��7uƖ7��O�!���Of�u�'�R��f�qO(���I�)+�Y� *C�}
|�)�i"�'剋!�l�O��'����S�,�� 2�&QguTdY��ˤj�����'ЂM����?��b���'�f��DO�	�M�(n�u���A*b7ͩ<���Ű{���'J��'���>y�o�?���ڴ"S?:~�\RG���]���?�5�E���'w�Q�H|�%@ȍ)��P�cv�0���`�����MK���?����A^�P�4ev�̹�D�bB���?h^)�ဘ�M�6����?IL>��_�'�?�Ǘ�;�Q2��S6���eΦw���'D"�'��]J�\�iUj����	;!�6-�>5��D�'����)�4|�O\y���?���O:���O�|H�a* Xj�`#�#Q_8�bl�ʦ����v%c�O<H�7O�D� !Z���5����;*��q�,�NŜ�*�BK��dR�w;��<Q���?������O�+��a��^>>��7��.Pi 4�f`�[}�,X��y�'���q����?	�$�\_B8��U"PV�h"��:]���M>���?Q����$�;O��y�'Df��Z�A�>�y��a��2���n���Iß`	'A���i�O�$QM����(��1(�)Z�Q����CF׫�T�'���'��V��@/Ӥ��'f� �8r�,�2���r��XHΰ$�i.b���~ҩV��4���D�O��*!�x㕍�#E������P�8]�7-�O����<��+�.�O����5f�L(.�����i�섩�DH�NHZ�	����k����O���?�i�M�u䓗)E��w:���Rksӌ�Qr��B�i�6�'�?1��^g�ɘ�JIs6�ӣ:P��(M�S�NQz���<Y��j����O�s���Y��Y�yc
�0��;{��p��r�������}��ޟd���?�(,O����Ob�qs!��]���Ƿq���K��n��q�d�ON��5��?�X8�#e��7Q46�ّ�ɷ`e�;׷i���'.be�61�剨[>���<�7`zӖP�lBY�捓"�T�G�z	e��z�'^�����O���0Xi����Mk�����N�O�tmZ���0�$�����$�'�L-)ɟ��ʣ�9#���0��֚(��z�#�I��'6��'��_���D�I3�`��D��V�F�� A�z��D�,O�Hk��'"������yZw��x�L�"]ę��
T��lz�4�?I>	����OXQ��H�?=H��$I���f�r�(yg,fӔ '�O��I�g��O�b\>�p�r�:�⠆�1��D��7�9�2�x�'_�IǟLk�B�g�t�'����^�K��y��ĄN��P��f���	1����m�W>A��N,�dK>ug�1�qHT��Rb͂n��&�'�	֟��F��z�$�'L���5�I1R���N	�Ty^�#��6#��	%(��$�ȭ�[��GxZw���7�!]�j$��� �UtI;�O��۠N٢��O��$�O�	�<Icb�	J�|y��4V��IQQn�@d4E����y�jX GxJ|�UBT�=�"0d_"4�i���٦iS3fӞ�M����?	���DZ�H��:�BAp+�8c�9#G��F�V���L��-SṼ������̖'��s����$e�j!��F�ԡg�$%���4�?����?it
A�I��	���O"���������h/O;o�m#��[�'ɼ�n�����{y��~��?����?qg#_2x"�),?´�hu�K����'D~��d)�<I�r>�	��@��O,�"��`۪%h�ʖ =b�i1�bӠ��?IJ>���?A*Oh˔-ܵUN
����+
�삂� ?lP�'� ���	6�X�CX>���Qr�ЀfL�E��%@�xF�pc�[�����uy�'��_� �ɞp��y��^��,�'�ܺԌ�q>؄lZ��h���<�@i���i�O>ʧI���o�
ww��UY$�J)(pAB�)�:Or���<���t���R,���č�����哟[قq���R:��q��i��O����'�哏1�On<��#ޑpvtA�4��-�2�¹i�2�'��I�o�b�詟&�d�O����WEz��`j�4�ؚ5i�XrrxIp4OtWǣ�?���^�1Dx��m��0��@�Y'(��7m�e�b��u�<˓ �i30�iYb�'&��O���O}Ac��1ʼ�rÃ�.~�T�%͘���ş ZDNh�'��9�A)�	�H�n�Ӑ
	q�	���0"��#�?W�T7��O��D�O����j���o���d��X�@4pu���(&�� S�N8Qʒl
KY��'u�	�E����|�����:fM�E���bǛL/Tl�E�i�"�'H�$\�G�6��O�T{� �O\�䊥_t��P	Bh�����1=$�$���LP�&�'}剭U���)��?y��BhT�BJ��0Z�{�'�U~� ���iZrW�6m�Oڴ�f�O���H�3��I򟛦O�AA��{���2&�{��N�����
����O����Oj�D�O����OV��6lU�@6a0W��93
>�"�ϷsZ��m�柀�f��t��^s����?�	ǟ�8g��=�:�+wD8y���0�[�|�t�I��������Iϟ��'n�SG>e���݆~0ё���ind���|Ө�s�3O0��O�>������$�O��r�]�lY��v�����d
T�^A��$�5�I��,�	���'{��k�~����1�QuJ��D�a{$�8�V榱���,�d��bVF��I��,j��e�h�'��\y��Ο[�|�Ó��#��,���p�4���O�6\��UW?������;���k"�ˡ0��%f*��(X�kqly��	�\�I,�R�Ia�	:�yW�*m���CL�"�Fiٶ�$�MK-O �zI��]��蟌���?iخOR� O�$��X�<�F,Um 	[Zf���O���g�ɞ*�O�]iP	<�h�ɀ��'}*�4{ĺi��)6wӸ�D�O������'���"�'5�,��HDH��[�Q"���,r�X,c7O8��<qĎ[Y�'�?��Nh2 � �Uq��ח�8���4�?����?�׍
'~�I�X�����O���D�i ���פ��i.z���M;2�B�(۴��%o�)�S��'��'�����6P� 1�%�,�h<��Il�T��s�B��'�b�͓�?��o�\c(����	�+��\���0�O��Ic��O���?���?i+O,��&.-\E���_�]�� ����%J����'��`��?2�{�d�'��BV:T����jH�Ez�'B��k�"5�P�'���ɟ��	����'��$��Cr>U�A��nH
(�z0 ��p��O^d�B�'�bƢ�~���?�-�.�0��a�H���_6��R�<ꮅEV���	Ɵ���hy"�j�������-��b��F.�w��1��o��!᩟��m�O����%!%,��?}��*x��<k�B�3�p��T�Y'�Mk��?�*O
Q�U�|�S���.xQfр�mǳV[�Q�bb(r�@�2�x�8˗C@����I����	r�I��y�<�P�K� �.<����J��M�*O&������mQ��������A�'J� ���-�4�*� j��<�\��*H�?Y��1�j�ً�B���'+N:u	@`T8erx�k@o���UnZ8#�X��4�?Q���?��'E��	���DS9(�3Ky�ܔ���a���nOrbM�	[�I�ʊc>��I�w��� ���	T��q��T�_�6��ܴ�?���?���C��ɡp
����O.��i���qA��
j;Z)$lŐ�Ժߴ��/����u����'B2�'l\�(�㍨+{���
�!y@"@�a�z��CT���'�e̓�?!r+�W�\c�TYc�Č��K�;=�N	H�O=�I�O�˓�?���?A/Oj�),���4c�������=Zo�͖'f�	���?���D��'�"�׶sH�٧n��eSG�j�����'��П���۟��'��5�'f{>mk�Nɀ}J��;BNH���O���'�� �~�'�?	�ʌ�{�uJX���@rX	��q9�\�|�	�����ay� δR$�������(/Bʹ:v�"r�:b�����}
�ɼ���|����	�����ŧ�;Vlĩ�uӈ�d�Orʓ :�T{�_?��I۟�ӽ���q�\�U��£��bK�EMk��A���t�IR�.�	ܟ��'�H�݅\U��7M�7-�&]*#/��O��6��<�D�����'\"�'��d,�>�b�Ռ\T��ckմO�&J�(R16BI����?!�A��<�����O(\|ȇH%C7�$K�k�X$P޴`IPP�R�i�B�'b�O��&��U̓��-h�+����IIX�¬z��H��M� �<Q�����:;u1���D�:㢜Aр�s�z<2�'��\m�ܟ��	ϟ̒�@����^;��D�OViAG�iEd};@*�phz�j�pN��b�O�
�������'1"�'�����_�z}x���/�މ�u&{����:	�(��'lJ[�'�r���y���5����<5��-FB �V��:���J�1OJ�$�O��$�<q�, /��V	�d*�v��}�-#'_�̰�)e�h��=����?	���D����]I"�¥F��*����]"�b�L��ʟ���hy��Р��g� ��O�*8�6�����>4�,7m���OV�
�9OD�)�O��О4 � <z�����,'xR�sw��2@�,��'��'�rQ�,��S����O���fG5u�p����C.���Vަ���*x��I�uD����Ο��%�7?��'��гpFԀ7�Xl�$@�)P�۴�?1���dP��8T�O�"�'��D�Z��b�N�5�Z`�t��tq �ɟ''�m�$�'��H@!�O�xͻJ��a�1�-k��dpC�Ouu��mZ~yBbP y�\6�O��$�O�IIK}��V�8�HA��:�4��!��l�F�'ab�P	�y����'t�K|2�P 1>��Q��C)ybJ�:�ئ�c��M����?I���WV��J4�O~ʶ`L�v=�������"q�Oئ��U)&?�(O�<�����O�<=#�O�1nܘ�E��e�q�4�?����?qDbקL-�I�q�����(�BMoӒ��D����tCr�����,ʗ�i��'��IW*�yʟ����O����i����	4�����ت3F��oџh�5_���DΠc�d�O||�p5O�������ʢ^ �T�݄7��r�_�h�O����˟��I����	[y��� 
��ytyP&kBLP�y����%Ϩ>�bkE�<���p�(�ϓ�*��?1������@Ɇ F��MC��ڑ�p`ϓ�?q��?9���?�(OhJE`]�|z�n�";}���M?:n�2�@�aiA�l�l�	)o��I�?=���x�2(�>!�
�v�\�W�\��H9pCM����͟�	㟬�'��=��@�~��Y8������q��J�bO�y=t��i�B���y"/ �2���'rr�{�'��R��Y�,�q,6����n�:m��� ��FyҠ����'�?���Rg�7EqJ(�TL�p���c�&p��̓KyN@���?y�Ɨ�<�L>3�XY�Œ�f�కi�$"ȸ��ij��'T���t�'=��';r�OE��ڒ�J�F�H=�g���)���q���&��t��;._e���V�	%N�$�R���&��0A�i�֑cr�i�����O@���>8�'�X�̧�X��3�R$f)��Y�� y��i.��r���O5h�1Ol�dG5�!,+�NQJb��+���o��Ж'<��P��'�덲�y��'i����4)�ԍ���p6l�aeϜ�_�h�����'�?	���?Y7.�V�a���A\�j�ގ1뛶�'dv�a��<��
r��	!B����m[�}J��S��](�%!�
|}b��Ҙ'��'��_��p�L!7,&����*E�@�8Q�Ń>j�i+Oĭ���'n�FJ��i�O��$"�\ Z�È2j��8����3�(�I&��O����O�ʓBj`��S7��ص)��-�E�G ��� �'M� ��?���@g?������	�Z(��S** ��j��!��oE<�A�'a�'zb�'r���0C�i*��' �9b$��Bu�D�T�./ƽw�i�N�DJ�f�*�ڵA����O��R��<��'�b��!���
�B7�R�h ���޴�?��?�7�d�8F�is��'�r�O?n�;�蘠�4��#��5\�Xx�QS-�R$(�yB�'K��ɟOB_�T�w�X�
U�Ƕ��� ;}R*��4�?i���	"��i/��'���O����'J�����vS�I�BY6'�4�p�*�#�y"�'@ y�F�$D���'��Q ��Z�'8;�b��\�Yܴ4�r�c��i���'��O��T�'�D�w�'/�� �B�����	�Uڙ��+i�<�j�%�<�*OZXӒ����8��]�!��k�l�<%�F���2�M����?����]�1�i��˔��'#�$1Y�� l!+��"\FVA����eܢ,������/1O����O��X�h�Јx�� �����D�:�n�؟��@.ۄ�M��t!< H���?p���|��禅�c�ï;ynl��區 ��8���>�#k�l~��'�R�'��'��\,Y��;`C]$��{�O�8�L㣯h�n��4�����O�q�;���9OX�dE�{�Ҁ�����Z�}I�)"�P�<I��?	���?���?)��@�%h�ih�傃�ޤO�mҕ-7P��T�c�z�&��Op���yP�D���$�O��*F8���G�� ;C���a�^a�E
ى�M#�'2�zY{g:��Z�]g,�=+�t(��8�RB�	�/(�XP%�X���q��{���ɷYĤ� 7��!�����gY
�:��|��H��iϵ[R~�iЦO)g�x�t��&�i��Ҷ(`���V��y���c���!7ؽ*A�B7[y�:���<6�Bɹ2ߠ8r��dݹwℵh��2d��)��h6���go�,F�$��@/�h�!P�D�#C�Rʃ�2���O��״g����N�,O���@�2P�4a�lw���1�̴���Ob�ܺ2�S���O�ĉ�%�!Ay�%���úh��ؒ�L/.p�c��כK����O?��@�s$L�g1k��AF��53��"�&�OB��8?%?�'�8��'~=D�sVoܥv��D?D�<��#֐#�j�j�5��c�;���<�� t����N~�+v�C��U��kȁHB�q���?y��[(L�������?)����$��|���P?	�4�ë�-k������m��dA۔I#�G6�T#Me�(�dɻ)�
��YȄ)RcM).:��ě�(�LTs�,F����h�d���D�G��d�O�el�?��?9.OZ1�ƣ�"-.h`��ɷtZ �aś��D{J|�>OT��kM�H�k�C��v^ꔓ�kԐ%�ޙm�i��n�Suyrf��s�x���T�a+�!v�Ę%�${�ʒ�=�"�'�"�'�D�{��^�b�?����A\��ep$Fئq�ʜ����� *d�qh��GX�퉘 :�����2m�&�� ��?�4!���8;�j�G��=9W��ğ �ɑY{@`1A���KZ��嬋	cp�E{R�	�W��Ql��CҤ|⑭ӏ
J#?���ӄ^dn{��]�{�jq0�CQ6�����Wyr��n"�iw�'�P>a�4�ْiE�@���A�Z{&Jf���$ɟh��4N֦\�@�y�!�C�L�w�ZM�S:Į ��]2<�����A�	�.A�8ʓ�R���K�.od��:ž�����2e��K�`�([W�
�`�´Ҥ�!�L������M3ži��Z>ux��/�MP$�S1T!��27Mş�	ß��	���SG�'^P1K� �\^��'Gۡ!c
a��'�$r��T?M)��Ď�M���D����c�Z͢pFJ�|p�x5F�0�B�ş��IY��݊b�'Kr�ĠY�@	)�6^
��e����㶮U <�!�N��)S�:���>�#�.4*�x`׏C�+�� ��2;��\���	�A�ɧ���BR�V~.)HEO̼{�d`1�g�5) ���'���'���Or@��IF�[�XxZA��D��)��4O@�D&�O�5b�I��E�,@ECXy��6�xbI}��(�N)��?�ji�T�1�ѿ%g�DD�ݳW�N�	ş8�0
����	�I�����萖ʝ�~^X ��y����VL�-=B��x�h���'�L�c#�fr�����zF{�%h�u�D,�\��2��m2��d��$ޘt3�
ّ
MDTI��hON0�RfϦR��9�AA/ �� ��O8��W�'nr�'3�OB˧e��X"%	�+��yr��V!��	��y�F ��X4Cԗe|����{������DM�~�V��+1ʞ�n�)��+b�5�%���X��@�]ӟ|��ϟ8�'Aı�#�'^�I�W/�t�tC]30=4�B�θ��` �Z¾L��1���Z1ǜ�:�JT�T�S0� �w��
`�Kv�4�O*8A�'�B5{:�tjs�J_��3�[MX��'��� �?�O^�a��kã$t$;k�=-�����${�O$<H�B*
zz|8�I���`lA�'I\I��'��IN|y]w|R�'��N�r����ݲ!f��,m�J�ď�r-���ៀ��
4{qP��3}���?)](�< ���Z6�n]��^|�'�(���.M�M��f��81��φ]�Q�`��/�O��$$���O0eA�"�8B	��*3�"���-�O��"~ΓG.T0�$Su�����/B�4�'��#=�OG��q�O�A�F���hʦ(��ER�&W�E)<Or�j���2v&�D�O"�'$9Xl����?���Ӫ�0�L��_��!�$ϺEl"����a�̋Ƃ֨@***��b���4_J(����	0Z0����`\@��mY|�6��C'N�00I�#؀^�X���O�D�0�v��x�	�/�X�C/�����O$�S�S͟��'ة��oȤR�>0(�+�/q@Z��'��y��D�)5��Y�(C�^U� HI<a�=OT	������I{��g��C��	�4�ߕ�
%���0x�FY�M���?	����C��Y�	�n��Fۭ��P%m�,K���������� � s�!�
�B�9SdR��*��O�d�W�'���x�jͺT�]����m����'lޭ����=�r"y؈f��	qT����w؟�;�'���0AN4\�x�j'��T��Qfc��O�T�9 �X3�Hم~�:�S�&�.v��Ȇ����a�F�/�3�jB�b�لȓ^HuE%4ʍ;�
�P���	�'���g��) J� �H�![6% �'�m��NA2OXP�f��?}.li�'�@��F�b	Tx�,P4@��%��'1B�
�H&
�����	6tm��'w�d�.7n�����贽
�'i�a)'
ܭuZ!q�-ܠ6q��'f�ES@�9�MK�m�"ND��''X�cu+;�F)���Lw� �'�z��%H�+;��uat��./U�<��'�,�2��|�z�,�<~���H�'���ʋ6}��ʡ�
�y����'}�aѣϸG�l�X���
B%P�
�'B�)�5$�}S�H!��7j�ҽ��'��l����<EpJ|��O�w�B��
�'v�*0�8���Q�Β�4���'��9��� �*T���Ц?պu
�'�z��=+N����K2�T�B�'�ޅ�Q�^nh�j#�O#'ׄ���'�b����8�܀��mڷ2��|b
�'4ĵ�A�A)\=�!��F!$D���'P�d��%��K @���[�>\�'��<##��s�:m��+ͩ��A�'�X��'�zT�DR���Y�TJ�'I��G�[R��@�I�J���'.v�Z�$/���z��VBμH�'��P �d�E����2����'��C'GL�{�,��,�)��`�'��sS ��q��S��dJ%{�'���;���E�)�P!�֮UH	�':�b׭��/ �cSϴz��	��'վ������p�u(�%J?=8��P�'�T��E 6��m�
C�@���'��k��`$y4	�>><�H3�'mz��ׄ
�)�0x#OZ5?���'��d�&���ɰ0Y$i�'��	 ��@#�o 9�2�I�'�y�A�Ё�
l���B)*�b�8�'TAh�ÙTA�qk�f
���K
�',u��l̄�>�P���Q����H�\�!<�S��t|P���F�z9X@���t�
���VK�L�g��r�zT��
"<����=���<	#H�5a�DT� JC#h�ѕJX(<Q$�	1jHٳ%9_���$IP	ff��P�'��)��D�10Lh�-ɛ)�X���(��p�}��\m� �!�߲T��y�����y�냀q�tH8�[2D��F����I�`� 9�?����7Uڰ2@�T�E�x@ö�n�<I�k-��J�Lɬ-�$˄��n���-|X���T#�\)�'똏7|Iƭ5$����IO�$SP� SB��XB��v[#��B≼#�4X�R�<k�T��׉�+\�B��>~P!c&nʿ���`�Y�
�xB�I�W�xhbbN3tn�e뚮��C�Is�F)cf��#4���"�M��xx�B�	o߫l��e�Ą<	v �
�'\�!s!�8o�I�I>1�!�Q��0���Qf��� ���	�$�OZ�U�>� ���GM�t�L�3O��Kg��RT"Ox� ��ޮa#8��p�N$}��4���I~���D���}0
!�!��D6Rpp -�y��@oQ����f�ͱ�d���D���㟢|r���k;��ǆS;���v�V�<�I�<�~�z�i]�O3�}A�jJ�I�K;�]��ɠ=�� Fh�>�9�A�m����٢5�����R�p�VՃ�i�`?`K�-:}K�2u@~� 
�Ql-bg+�l3��7�[��QD2���Lg�N(�`w`��3r%ۑ�F�w-��%��/6�9g
O����� ] ��T�\eRX��Q�``�Mt~�>\�X�D��,'�O�>����ۍt-����.7�*�'����сY+��0�0GS"�8��'����V��H�$�c�)�>�O�H
Ô?mA�
�](�k�C�4�`��(�O�LD
'�
��a�,�q��A<fAs��O�a3p�ˤT8�	�5�?#<1&
���-1�3I��pX-�G����ȓ��	{D�üt�8u���*6��!D���<�Is�'���@eW8H ��O bo`����+ ��DmG?Q�H��_ "��S&:ǘ�ؠ������J�6I��B�IUJ��qO�3-����9���R�� 8[w�=a��Z�n�����O�|��O�1%���8���V�l�U��G� Qg��~	�C�	�	7��Ԟ;d���Q�?!v��t�a�ް�w�\�w����#̞�|2����?9��8}���Rn@g��l a���0>�dc*UL��wo���u�C_tRɘP�:-Rxxd#L�}��43�/���?�S"$���z���O��a4<_�������!\�)i���emf�s+�((��}k7	�Oø�������)�o5DM��B�y!b�[��M�RY�N��:7	s�ax�S�d��|��o]�z[����-Q%�0�	�fܵ>}�4����9[YT��Ӻs�_�q�������4�ˑ��h�a��B�r91� O�L�Bm� g�f5��`R���*��4oT��ɎF3m(��@0�p��'�v��ʒC?�ݻ:$2Z'�ҁ� �&w椰�
�@p4�1#�ݴ7�t)v�־fu@ ����#MTTu��� n�O���	_#�yҤ( ���=Q� -_b1�IXwm��򃡚a�'�0U1��.>�`r��Pn�I��Ӻ+ �B���HRBq mcF��g��`T�~��#�&��z"I
�<_��B�,��O6�T'�P�5�a���TH�X�`kY�0
4Y��|�X:��Y�`��-�I��i��D%B�z#A�p=�'A�7^�J�O��v�X�er���T&V��,q�B^�!g��S�4P����ļeNZ��|� �<�;Eq�ibc�POx�11�	�z-���<15��:���P�.�xd�JҢ�1$^ݓ���;n�k�O���~�⎜	��3+OZ��2���&�{O��`3�F�/�����$^�T���q�+v�l��F��13_��)���@�Ρ2En��kO �VmV/ȼEo@�0�Xi�'C@�T���+r�D�*�p<A�	�E��,�q=B��׆K�	!1�B��ӎ+$��6H�AH1O��H��!��P�Pĕ�FD�Ȥ��,W����I1�x�*��Z3�$��s&��`�2	��x�Báz�(;c�Ϧ=��&�_�S�t׋W�ԑ�wIvU��C�qwess�-A�S�yr���Q�lGe�'�$)V�A*P��xҷ�S7�(J�>�(O��w(Y�Z�R��ϓ�-�0��]�t�j�I�$;e�V�~�6�3Y�| `���ɲ$',Ԩҧ� ��I�&Q���g.�B,b`�W˂(.8�Tk�H=f�1(�*�?5,����ZU�'���1I=Jw�uc5�28�X�8I>a1�xtX�:��:��?�HeEF�LE�gBơ M�hS�B��dUEM�)Y5+f�]q?�"���!2����+Vt�J�g�n2]"�)"�G"|�杊6f1���\d�M@��5*b�LB��5W�*��d�Ɍ/�F4K�O=CRn���"Y+v{�4�O�˓}�|�0�I�o���rcԴUIZ��'��Ԯܞ`@��[�
^
I�#��m�O��'��d
%�.�*y+�O��1�i�1K�@�2wiÌ
� xҧ�Y>F�pD36ͪ��=ʘ�?6�2X�Tq�B^Up`]Тo+!S�I*9�T��qI��,��g��?�0E�ӝB�X@q�,���D:2DV-t<܇�	�@�z�a��0�y�ˑ($�>��"J99m^�t�%f8�@v�3ғ���Ŋ��Y`�w&��DH��0 ����{Q���}�N�Cfh�:��A�3?�	M�@D��)L���I��by�HPy���!�e@��A�4iȻ��$�r�ؤ�נ�3�c��L��q8T(Ǩ�z6MȲ0�|7-�C�d��<��jH��
�A�l{ DF�.�0#���aJ����ږG�d��6�q�axBG�9t�	�IB�6�!'+��Z�TQ
M�l��������T6͕�P�D)ꌺzwh���#λ71\�		ϓ:�h���+ޛw�GG�	J�J���b�$���i�@��^�r��>��O뎥��Is��"%�z�g��E�? ��r�<n���S��e"����d�(/�� X$�4s�H!�^5��'�*Yi��՛��Y���3J�h1�����X���ů�P�H>�;+@�qJ�ɦg�Z
�h4,P9dB�ɹ�a��,�ܣ��A�C�A"�����<�*�;uה�0DF�Du�`)�I_����a+�A/O��y�c�iS0��L�N�"���{x�0��D�/)"��6OH8� ��T�!;��Öb=2�0�����<9��Ӷ"�2�2��w��̻Q�O�6uv�[�j��CExZ���ҁb<��2lέ���b��u^]K��#2�Zi8�/�tߨb��Id�j��xSp%�/l��h��0���
���
&�P�6"d���pVTۈ 2��;��Uډ��j8}���q�,�8���C{�6o	�h����R�cY�83�/̩)s����)*9,��c��2w� ��$�%$� �O ��,��p<�e"F��}(ǶO���ō���yזS��͝�<�%V+�3&�ߑ^��G��!o�b��ϱ �C����e+�"A\��@Q'�-E�rMv��{ܓ9&���M�W�2˓
�'`ֽ��F�*"c�q��� 8f��z�}"�9/(^�[�f[;5*���å��� �z��1a.F��	F�6��lV�_����'UړO�)b��$��$���>-��%]-`xI&AX�\��aԊ	<����F�'�jD��J+<�; ���|�}��6�DP#Sy<��ǓQ�YP�H��d�@�Z;x��8�`�%E4�1a�O��HO�|"f���I!=���Bm�x۶Pq��[����'����`Z��fD�V��P`FE�jv,�J�aB
��'�<MJ%Θ�K,�I{n�'Y�U����c�����E*~�D�Ҏ���hU:d"�n��Gl�z�*�9"ph�֥B�[{v�����4��@AϗMS>H��o�-���'�6L�L���Ĉ J��q�L=3�@ޤ7�L5�m��%wʼ��'��l8��D�]�IYv��1<L<1�H΄��'��h"ႮOK��
�Nq�$��Qn�:K��K�G��]qNۆ*��%�'�&y��!qpB�Qg�l���M@�'���K�A�6���V�s��kR��4Ue 0����$k�l4:��3��$_^0+p"۫@�*Y`*Ѐ��'�X�0h�&��˓ *O�!2g�ч<9@��@��':17�'6�:Ձ�ae���/͂t�H��FCȩ ׄX�W��e�-Js�T?�?	tE�e�Z�N�>]8 ̜�T�胱��>�"�3ej3�5&Ll�t�)0��kM�=��D��?ӐG"1��y���Y���Ǥ0�Ɍ=
�Ņ�	",׼��$,�|󚐁�,A% C!�v��BBA�3�9LU 4l�OQ>睈f��Q0"K�,a��h�a�Z�zH�B�IT�,p�L�<���c���$�BQ��O��B�Y~1�Ab>r��IOH�Lg�xd�c������$[=;����a(�dȆ�H��	X
�`�F�q�����nجT.n����.�p>�����&�w�0i@�x�'��a�'F�K���3Dwn^b�S���0�$]�F�)l���)j�<o
g,Z�<[�lh�d�#2)^��3�V�X����V�fφ< ���OQ>�+N�$	ej�_=^���ԪlD�C�	�lq�����Ȑ�XFN�f�Q��?��k���!T�%)eN�?�GzbD,n��Y��҆#�@}@�ɻ�y�m�+�X�@N�	�>�ڧ���y"O_.w�LԘ劉�U� ��k3�y�H���!�)S+x҆oE��y�'C(H�=E@ǃM$<[sԵ�y�S�c�
�hn@�M�fy��Fư�y�H��\��ܷAU(�s���y�*_��Z("��9F����Mޅ�y⦃/�^4�����#
!*�.�&�y�^�X0�IxG^-
��@7�#�y�a	U�pp��U�{�2��W �$�y
�,]nN	�"#E�AO�r�\�y��0o���Uj��;���#��Ӭ�yb�יb�5c��:\y2�e�yB��<H<dIP�Ŗ2�ZX��J��y2�P�>c�t�o�4+���qU�5�y���� �:3G��W�P� uG���y�*U�BS�i�aN�%��#c��yr@ͼ����!̇�0��%Z����yr��"�x}*S�8<� "�P	�ybM����X��I2:FTl� b�yB�s���2���'5
uZ3J���y
� 0���ܮ�Rm�CjT>E�"O�5��'ʄf ����`ֳeQ�M*�"O �C���]1t�q�hPm�E�"O��+�!;��)��4|fΔB�"O�TrQb_5���	'b]�� "OQ�/F�	Y~]p�HH�%AZ��"O��sD�4P�ŲW�E���Ѱ"O���ğo��8�'�Q- o�ȳ�"O��t��Jo�����>}�0�p�"O�,Z����{"����r�|�V"O.y����!>j�;��I%"t��"O�؉�NV�*7L*An��b�h`�"Oj�z���z��|��*ջ(����S"O*X0�٢E#V�91h^�k�$�9�"O�ܘ�e�2����G�,����"O\l�w�"�FIDF��P�Ԡs"OF,2pHԩ'�=�����ng&�kt"O�%�c�j)k�cX2,���"OVm:"&��}���ڂs���"Ol���R��fU�E�J�Q�"O��IP�>Оj�L<H?P��@"Oά8c�;~L|a�Ԣ.,<)�s"Obx��B'i��}��*��@���"O��-ZC��`;q��D�h��3"O:GN/[�!��c@�k��Kq"Od�#�C�T��a�P��	1�jP��"O EY`hD<;~�9�n��H��"O�������2,����\<�%"O�y���$P]n�K ��=�H�"OZ�ӓF���<Z� ���qC"O�D��D50��d��iߒ��t�"O^� �Z
~:���VCĈ.��Ȉ�"Op�AĢ�<�Ī�k�����"O(��-ͱ�����`��#E��"O�s�j�M�Ԉ��@�b+}3`"OD���P2��1�]�%Kn��T"O�=� �^s��A�;'а�"On!i�,ߓ�f�:���)*f���4"OK�!�4���MاP���L	�y��Y	o�� �>q�xqH���yb�NK�v�z�$Z�U����ԟ�yb���w~��;t���x�CD��yR��O&P0�"Iٶ}Z2Ȃs�ڛ�y�#��|�x�C�Ã�u��D#gҚ�y"�2t)V�'Y�p),4)Co��y�Gn$'�^��9Rׯ�4�yBgÃ�>|!�e#X B��BF!�d�,a����7�iI��Z>3!�+l���D�T
�B�@�!�D/���2h>$������ِJ!�$��	��
SR�
���ct�ӧ!!�$ہx��ԙ#�2u�.09�,(u�!�D]/k�jb�å�L�#��$^���Ă���3�9A�����דg�8C�I9o�H�Íž+d�3.Z/0�4C�I :}�%IF�<Y&i2���l?C�*Iv\8R&��+a��������D�.h�f�(�-�8/�lP�`͑+�!�Ϲi�$���a�n@2x����3�!�D�L�B�tg߇D��Õ��+m�!�DS��	0�d��H�L �!d��]�!�D݇,B	�t�c����!��X.p^��A��?���[�gI�!�B;)�\�s������F݉o !�� �q	��ӣ.FP$�B�KR-� "O��Kp��-u�HV��%Eи��"O��#��T�P�����Y# K�@��"O�\�j�,Fij J��g1��k�"OAB��,�*�Q%�	\*pD"�"O�S�c[�0��B�E��`&��R
�'��j��(�~� � W����:
�'_*X�`��C�^\ڄ�ɻ~���Y	�'�<�8�&�o�h4��iU�gb��C�'�~��Ei[8b��I�Q"^� ���'Cʰ9�&T0K��0�L�b�D�R�'p6�H1b�:mf�8'��6]غ�+�'��1	C�N$S�iyF"�Tx���
�'���Dc�5��ًe�փY�и[
�'JrKEI�" ��4�ȜB�S�'�:�f؍~KD��P 6�����'�ZԺ@N<��ٰ�e?vh	��'�fd��,Ƅ&Y��k b��$!���'�(�Y�7p�}Bs	F�h���a�'P��y�'ş�8,zU��7n�4���')�##G��~pXJ��P_hh a��D),O���E䟠D�=�����k�l��"O�q�gf\�W~��Pl�W���T"O$�Cqȓ�Ha�� �d�G"O�4�Ko-�P���W�$��C"O�=9��84 ֩���Q�~�0�"O��rd���*
8Ms�O�=J��Ń�"OP5j��V8$`���f�ߖ\0Z�k�>ي��i��<u�-�eH/�`�i C��!�$Q�Je�AKF�$��؀���q�!�D@�G��P�%eP1Ux���#��!��ٙE�،�Æ2�N �g ҹF�!���6Iޮ5��V��������d�!�$<8�vq��C�I��ɋ7IJ�m�!��hȬ�3/�����eʘ��!�$G�K��x�,��f|���V�|�!�좨P4"�%n��ʗ�W/[�!�D��z\B�BZ4TQv�8�+Q<Y�!�Ā5%;������ʼ)ꌬJ�!��C�4��@��B�p�r�b�Q�Z�qOH��䝝0S��&��<���g�*�!�䝚b4����՗�6�#��I�z�!�X�us<�/���̪o@��!��M���9���@������O�!��C�E�����Z�,���cjD��!�+wJ�S�Z���e����)8�!�$�^x���b�:1誩��C�-�!���|�,�i5*�5V��A��\�!�DO�P�N�Yc	�Ԉc���!�!�	6A���V�(i#ЯƦJA!�d�9�FD0�%�;*�1
Я_�7,!�d>���,i(J�1�Й-�!�$}�H���Q3!-��j��ݠV!�dS�c �Cf���N>X�쟂=�!�Ċ`� ``P��1ې���(	�!�d�)�T�p&h� �6a�k�R�!�ןF$;�2��Iㆨ(�!򤑇]���J�+�H����a��Y�!��'�TdrW[�s�F�Ce@2��z����8 �a� ]�<�ԙY��6�!�$U0��Y��"����O���!�DL�	�|h{#%��Q���7`!��Ң������X��;�!O�T�!���T���,JG�8}��-�+q�!�� z1���բEOx�맬5M�0U�b"Odp�7EGH�`H��J��9 ص80"O`h�����p��Z; �pHU"O��@�A6N�``�J]�8����E"Oe2�gN�m0���	�
^�p��"O��@��R�-�r��`I�1+��S�"OFͱ2i��~�,q#��MI�`�2"O��6�ۮ?�6�(���J��5R$"O�%���b+���,��H�
3"O�(�`�z��I�TX�����"O�� @�ϑv�(\֊Q�A{�A��"O��P���g��D�L?bFp�@"O��i؃G��`�B}��o��y�b��N�����c8?$����
ϰ�yR�Z�z�2I"6M��0/ʸ������y���R$��jR$I+<�R�K�Z��yb���m�ұM�<3�ЅkUB��y�F�qAN��3�ǿ)i`-���/���hO��2fiL�@�-�1��9-,�����F�d(]�#�E���u06#�yR�R�d��9�t�ӫi��φ�y��N$�0\���)���U�y�@�pq�i@����E޾�yr/Ǒ:���b�1'D���9�y�n]=y��+S��LWz�#�ʓ�y�dB�/d\#K�3X���`l���y�N��|P�%&U�e��1링�~��'>��"��/�lQ榕�,h�3�'�a��K��s��vazh��'��)�g��dq�צ���Tph�'��9�wOF�62�u�v%�9~�L�z�'
�Ⱟ�`a�B݄@@�'+�����TaC�'��.�R�'y�"h��v����LyI�U��'3��q�⑧�0;Am$:�|�"�'5V���A�P�<���Z�c�B���'8(Y��A�$`�QBg�Ԩ`b� ��'���##�؎Y к'��!X�$��'f�|�p�U#9�6 �wn�V�x����#,O���l[�<́҅LieY*�AU�<�с_B��X��,B�qp1f�P�<!f"�\�!FO�2�yKsa�h�<��e a�~=KC�I�Ve��!$�e�<i�N��U�z�bc�|�JDi�<��ۘ/��)֪��H��]�B�e�<��M=P	����V�cv6EyQK�c�<�6)��"v�����q����z�<9%H#~ZjU���LTMZ0����s�<�b$ň^�<��b���`P��H�<y�(�N�,�FŇ~��-0��O�<���'1L�`�'�?O*ʘ��I�<�vb�m��\B��F7D�P��H�<��ִ�0����&��!����A�<A�A�)�B<���P%%Nd%���W�<� ��RW��1|� c4�,��B�>���K�Ʌ(s��h�QjtB�9R�8�h��I�BX4-9��D��jB�ɠU�KMjQ��j��\ ]رʒ"O���n2`�nu�S��U	���"OJ<rWM�)ߨd�D쉿{�����"O��X���/���Q��"a�� e"Oz�5�O�_���#g)�'=�h�"OVM#Ā0(�@hC��A�"Odq� ʋHz2�f'�$J ��"O� ���3��K� $f���\E�&"OP�RsN�L�$��W�J,|�B`�"O4�Xǥ��s����d�}TDtXC"O�A�NNX�!HQ�a.Y[�"O4T�B��6Td�e`�`O�jx�l�%"O�۠*PQ���	P@L�bf��"O�Q0����Kbm�b�?^L2�# "Oԁ8߾�*��V`F�&B	�u"OR��I�()m��P��A�@�"O��30n]7~v�|�B�,%$��"O��W�p)ᎈb���ƛ
?_!��8|�dPj��ҮC�^ܠ'䚰�!򄃝}�@�	@��)����!��Y�j��e/*L�J}���V-!�$f&��2TUEz(��C�L!���K�!z�^Q:��bM�!��	�J�
���Q�U���#�gNz�!�d�2�659���/�� $e	f�!�C�L�
2�H�e�PH��Q�j�!���%f>���E�XĬ���C$�!�Dȿ>�B`zv�(q�B�[?{!�ۄ*B�0 ��h���pEC�#l!��ÈQ<p�)e�\�`Wl7�!��?p뾍2��Y%3�T�;��� �!�Dǖ_�����B4Ѯ5���/g�!�$>O�ru�-��j�|�c�Ԡh�!��\ ��}��-�8��Bm�!�B87��� �41�]
%�W�G�!��6��M�wO��'"Ҧ悃k�!��k�MRL�(��N��M�!�d�'��E�wJ��\U{w.��a!�_#8�>�2e�$��RBM\�I!��>h��{�`-�h,�KQ�1!�DΊ��5rL0V��L���	��!�d�,��1A�Ig���(^��!�D�
����,����� !�dF�!�%��!T"f�����A�J!�D�t�A�a-�?�24���N=L�!��Z�,��$�`�Amp���&�3�!�5~�����*���R�&�-:�!��S���Xġ�/��i�2�_lB�� 3v����%�.��l�eh>�xC�ɵPzyX%hB�z1��k�HYbC��ڌ��JZ$\���5�ŝ+B0C�ɣ=��TX2'0Q���Z��B�	�Z�����AC�8bACZhC䉚!n�+�Nn��qq���\�&C�	�e�.���\�0� IF쇖+�<B�KSlC�M��)���J�D�;���Ka�ڴHG'�MF`"��W!�d�����T���|B8Ȱ�ڌ6�!�d�n\~-
v�3l,�#O7}�!�dU�O���0�̄Ok�Isc��>K!�ď=���!(+`ix3D,�41!�D�3U$4�6-��dM�e�P��N�!��aɾ���22ڼ@ToZ�!��=|��Q�f��<b2�x#@�:0�!�$�6{�
pK7AZ�~h@�n|�!��N�?:=2�koL�����.@!��Zpu�!̏jr�D��Q5!���'y������;fF��S:!��{T<x2���$�H�"ĀL�!�ſK\�		��Ҟr���"a��3\�!�R H4�c&G9Q��qPaS `Z!�� l�ɠME.�N� 0���~��8�"Ov<�!oQ�dB,�ujN!�8�"O�mc@+ų�b!�rlճk�p�Z"O*I�&�l�2H��-�An!PW"O�#�����m3`� �k "O��7'U8_�����
C���S "O��BbW�Hed9ˡjT�F�(���"O�����K/hJ��be�W�,���1b"O���@��l�|q֮��uՖ�+b"OR�)VOQ?A����I*v�ʭ�Q"O$ �g�]��y:!l�t�x�1�*O$���ޠwp�u˛�{e�Y�'
��ڲ��-Y�A(эǅxt��#�'���$Nbf�h�b� }`+�'A�uA���$r��|a��\4u�&@��'+��p�G�*F�A����mx�K
�'�<u�.��{B�3Ԭ۲UL�:�'���@�ͰV^���#�U-�T��'�P9��cZ/P5|P��Nȑ���'�]c�+�  �>h�@#Q
�>���'h(EHu��B�~Qc�E\�}PRD��'����W''�\<��G
%?l���'p��`E���P�D�B1T�̐�'� (�0�I�~(V���`O�%���'��ksK��=����m2gt�(�'��"VI>h�*ѶZ|@�Q�'�ZD2@b}h���]�Zup�'�h���̥ȶ����'2��X	�'���5���gI<-�������'�j�3��H��X�pmʻv�tt��'� ���"X�z���B�苾m�< ��'?2)��� P�����R�mr�!�'՚k��;WT��aEO!t�� b�'� cƇPy �0��ۏe��q
�'�jm��ۉ]�0�Х��X�l	�'l>1���1H�LH)!U�,�Q	�'t�E�v, #��` ZS���1�'��僥���p�� ��*<����'�J%z��F�aH�d)(�@ �'HtE9�Ȁ�z�,�1iW��6�8�'Ì0Ɂ���Zb���O���|���'Z�50�U�-��	�2��W�.d��'8��"C�Y="p����C��p��'��2���6(J�)��×�cpt��'gVl���20���҄ �_��9�
�'Ft���(�����ǫY�*��	�'r�HGo^�v,UK�E�?	J�`��'`�0P6"ʃyP"��B��K:6���'p�`��W�\�,I'F	�?t0Y��' ���$ֈ[�^-� �1��X�'_����W%o�I��(@�]�x
�'_lL:�N3K1�£K�]��
�'� VɊv��� 1�ϵD���r	�'�����M�O<4��0�Ʌ5��5��'*�a��B�O��@�`�.1DX��
�'����t��.8��S�#ފ<�.I�	�'$�2@f� �N�@bg׭.�2�'���cԤH>U"�B�$ T�1�
�'�rHI���tM9p!g���\�q
�'L8U�%����q� oȎ|���
�'��<��U��Xk�[
��	�'��t�WH@#㔈���+��)S	�'˂���eH&�SJ$�r�	�']�8�B��Ҩ��lY%	ErI*��� �`�6�̪C�=��/�&s�r�b�"O��Jf�1R��i�W6��"O
m3��
[��Y�9�$�"O
M;f�2Mz]	���M����"Ol�
eN�&��D�� �6%�G"OxQI����C��	�"g6~�*y��"OZ,����f�ش�g9P�ib�"O�{�æc\�����7y�Uc�"O�i�țB��)*��T6vK��"O�I�q��>NdYPN+3/$|c�"O��
�N�;v|2�͆�m��#t"O�}ɓK���#Z*��+�"O�9qТ�%%)xa3Bj��d�#"O�\0�d#c2�VA�9�|�""Ov���P6Ҹ�u���#�0#�"O�t��#ْ��h�ȣ9�N�R@"O��[�*TPG�� �h("O
8��B�$�%���<'�na)"Or���#�	E����Cәq�|�x�"O��е	R�7��9��1Cnp8"O��FM'Ny~ "@�Y�[Ɍ��"OPX[��A+Pt�ɳ�O͸8t��"O
��d`	'v���/�n�2�c"O�A*"h��AN>�6����I�"O�m�Β�H\k��X�{�x�Iq"Or�1��:!��VK*�^��"OF�J�`" d :���.h��V"O��q��1w����+�ň���z�����釡#W�:3�_%JQ�U��)�)�y�%�	Y�4���%Z�E�(G��y"�N�fF��#�IN�0�.S�yb�̧2	J����SDF8*��y�e��N�%��2}p�U)ں��'�az��RaW� !E@��Y���ϒ�y��9���[��%M��I�§���hO��A��0dRN��4�RQr�0�ԨÔ���1�O���& %iJ��)a	�z��@"O�p)���9>�0��b����"Ob�
`L`�2�hm͓�T��"O(0��L�@�~EBS뒹aۀ��S�|��'�az��Z��Qʐ�A��m�5���y����H�Q�ڪ�R�!��y���S�P��
�1z���C�)��d(�Onq(�ɛ<&�:+���pg�:�"O�T��L�8��Mp�(�$�>�b�"O̤�Մ�6ފ99�?��1E"On�*�����L�B%u3�`h��$LO"�82fP�cZ�@�]C�4��"OJ�{0�E�Wm��G -���pO��f��f�Д5��$�5pS�)D�@��Q3CNP�c/D��-�E�4����h��I�� @�"@�,�tYGo ��C�����/�1sf�0Pk�'��s�'[�����rKD�� ۗ$�@|���x��06 1�"A�+w#R����y���G���{�Y�lF��O���xR��y8��R��V,r�~�/��!�DX~ Z��Ac�5L�����%j)���*�g?�r�ݩ%���H��U�lf����H�<�u�APz|i��[/��܃�Rk�<i5A�DiV���rj��*�P�<Y#@*���ЌWXg�;d�T�'3ax��a�d=��P�v��u�%�ȱ�y҂�:k�"��dY�}b9��ۉ�?a��� ��+�a� N�yt��8�j=�"O^'J��V} 1R�)��4"O,q	��T�09f5�v����m �"O�	��iX;|��.I�?�B��"O6#@c��) 0�	fN�61�����"O�� ��n�}��,F�j�� �3"O*SN�xh�	��ĹF�Q�t"O����M0\�.��a�� �2U@��'�ў"~�B�U��Y�d-R�(*�e�'�y��X�6�z��EَM�@��:�y.�k0�H�j�7H��j��@��y",Ӣ~~H���UJ�|(�EC.�y���V:���a"�O����ĈG��yb�!a�X��pOJ�GV\�����?���0F�vm�5N2}� ��_�̰��?���0<	$��'It�R�F_6�H�e�I�<�1%�6f�$lCB�<E�ApC�[z�<�ޅ>f��m���m!b�FB�':?mkЪ�L�h��#F,��|q/$D���3(�#X$�4�Fo�	�bL �%|O�$-?���9s��=��@�s���h�OL�'axrEC�c�����X2D���'[>Q�C�ޥI�ba0pF�7��'�>샆*a���"nB~���5"Oz�S��p�0�0q�ġO�����Q>i&�+�@�[�)�s�����O��)�I^�'m2�瓑[Є�ŠH#0������=I�Od��~.�C���G���	Q�O�6l9��~{�za��/�.��'G�` �H ��s�N��Qo����'Q�4�E$�G,��
[�
@<:�'�0�±dʷ.1x�b�j֝*o ���d#O�,T�R�P!��L��(�e��(�ynٙ�Mi�?L��h��J0��'��O�c��� #�]FL8I�G�h���Ĉ.D�y���7.��F�s@����,D����J��D�i:�Ξ�L8��c.D��V��(��\�2%�� S@�;�$?D��Cֆϑ{XC�=����i*D��+� �4E��xi����$'$D���1!�!/Y��k͌``�Tg%D�\�vo@0t�w�I)6F���f,�<Y���S?"���K��Le*d���N�"�RC䉓KU�QD)u�V4���C�I�B�p�$�/.��L�TFچ:�C���q�v�Vky���t�۴Y�B�I�S�|�q˝81�B�Y F�2Ry�B�5�>��w���	��`�t�*F��C�I9PX����PU�r���C�~��C�I4 ojM
���9�4u��� �C�	.:Ya��Q�]�9!�	R�PC�ɐBɼ�@7c�r&�0�d	8	�`C�)Y��{�J�5��$J�+ȣrt:��$� ��P��+���h�3c�6D�P��N�J���z�o^<X`(�)D����`�,Sb���pg�pi*q�&D�dj@-K�(-��$�n�"��G$D�H�U����R�b�؆jH�#D�8X�N(��	�R�4K��XU !D�y��ZX�p�e �p�@)D��
_4^��5����1SZ���=D�����	4r΁ж��&4
�Se:D�l�@Ŗ�<X�3/��L���T	:D���+\�}wڤQa�Bb�*��CB-D�� ~��U�[�{�v�:�B�1�b�(d"Oa��+�<��u�[��m��"OQ�r�X�TZ�#	�B�.��	�'>��)T�[ր0(��1SA��1�'�Y�h�I��32,� :[�t��'Ku(���2ь�!���7��"�'b4��$OS�~�y��a�?��'w�\�0��,������4~�9��'��ܲ3)_I����u�WN���'xTR+�>�`��E!�B�J�2�)��ˊ Gnٛg����������0>��mO=L��|C�*��r�T󷁇[�<�D�ؕ��i�ő��"soW�<�#�pa�(a /�B鼝
�lOW�<A�Kε z(�ƥ�`&24/�R�<a��H<�̤`ǃ�k��"�RN�<a&	�-�(��VD
>����\A��hO�'qώd0�\�c�H�*���m�:\�ȓC�0PF$��b�,1�UA�au�Ȅȓ�0��#R!"	*	��	�e�����d� D���аk�*@���q�舉"A�
ss){v�E	�ZL�ȓhz0�;�o[;Lc�ޔBxࠄȓ}:��G2P��8�(J�w�m��Z����N��i�(�jfR7֚�
(O����I��N�8���E�P��b�M/�!�䖓FD�d0�]�S����)B�!�D�,f��D;�d\W���Bs Z�!򤊺-~�XF�P8`s���4O!�$��!T�{E�[�pd�4fK!�d��	/�� c !�:a��	1!��<B�`�2g�
�<�3 �#!�d��.�`Pc���U�6���	�6!��L?��pԬ޳aB-0է~!��Vn��pQ��6M>A��F�*!�dR�����K[
8��ꤨ�e!�ęIZM���
Q��@&b��z�!�;!�.و�"I'W8�����,3!�d]
HE�[��]/ ��ۂ��T%!�D�&S�4a��ڊS��A��߷o!�yi �S祕:L<�@*�=	���	..����E��Br\{bË9f�C�	1&P�,j��Z=��X��^6(��C��:�p�jW���v���O�2͚C�ɅU�)���5^���c!L�.��C��	�2,���ط^���C�b B�Ɇc�R���O�i��`���Rz�C䉱�e���!^����s�B�s�B�	�Z�
Xsԩ	Mk�@b�#1i2,C�6X�a�5�HZ��zI��U]�B�	+I��+q�֞L^�IvF��NB䉇t*����K<KM�p�D�U .B�	^�<�5���5��@PeEN^��C�ɅF����'2�h�0��5"�B�Ig��@�H֡f2<� �F�;�C��>a�*�Ȑ���P�+�"�ttC�<�քe-�k���S�H(B2>C�; Ԋ3%��^�`9*F!

C�ɘK
�5���ț�,E�YTхȓ	������I	���T�T�]9���ȓa�$xS#'�MA\���O`�Մȓ-���ٻ��hU���Ff��	P�����t�W�?e����D�_5DX2�:�'D���S��17��a0��!�DoȝN;!�� �� �VB��щ�
"�̈��"O��+���(
�&��-�$W���1q"O��)��5|i�u�M'F̜(��"O�,c!ɌC�v%;wn�
�T�Qg"O8�ڌ6ʲX2O�'5w�4"O��"��J�0���C�UBe�"O�!��&x]`Cm�h��"O|	��E� �����0j��i�"O(��,�-\@���9f�
���'��$(�`�����n�H@�A`�:�!��?X9���D��	.\����P�Y�!����|Xs�E=�AT� b�!�d��4��H�7n�
�(����!���!oA���p��t�r�T�п�!�D�1Y��0�NS?-��%b2�*y�!�d_7��	�H/�� J��"���>Or�� 1-�����;;� 	E"O�i�FZ�٠t�DJ�N$ �"OZ �2�ݼw��6F���ҘD"O�`���$B؎���
�*�f�b�"ODѣ�J�hx�,80 Ɏ+q<H��"OjS�"#g�}��r�V�T"O�Y���%=�	�E�'��育"O�j��ܤ8�jt�%�F�hv��"O�}���2Ѯ]�EF/3[��"Oc�i�4"<�q�	�O+�<��"O�t꒭K�7I���iǔAt�a��"O��QF�)0�t�cfȗl�y��"O��!҅N{���CZ u_|��C"O^���6���s�ʎEo@���"O0:�[���[���c�����"O����NH�%B4��V�k�|HK�"O�=`�T�\*� 4#B� �)���	J�DXP�'[��(g�O";��Q��"D�īf@�Z�0���N�9���C�� D�1�+��L�~PH����02�!D��I@	@/r2�ѹ���1:1f5�n%D�H�qa�%�Q����/j?�P24�>D������
8I'	Q�q�b���<D��<uLQH�-̮C�x��D:��n��@�3#ܜ>����󄏟�$�H� 8D�p��"�S*��0Ѿ𱀲e5D�TYdć�=�>S��� 4�)@�d'D����Ͻ��)V�LR�tA��&D���'��B��Z���/6f`q�"D�@[I\I=�8R�i�cE<X�� �D%�O.��ΖOZ�+��0W�p�"OF����aQ"�aP�Q?8-�QA"O��2a��pı瀝R��Qc"O*�1%��>�0����sj;"O��0&^��R�0��H�cO�Tab"O��E3[��B��;F(|��"OdX+�S�*�A�rf�(ҩ[�"OQy�J��S`yb�+eP93"O��;Շ�P��׀U����A"O~	�Če�\�/¿B�"���"O�)��eG�F��|:�Ǹ*s
�q&"OF�+t��� �;L� BFZh�"Od\���"o�B��B�0/B�5�u"O
�ӢQ�ii~ب�j"��4""O�D�7�� ^�����^�Ucp��u"O���'�K�P�,,��B	�:_��A"O��"o�K'eX�*FK:D˄"O�I�ǏC�?(�&*��F�p��"O� �Q�6��~0�p#�c�<6�.�c�"O� ٤�\6l�J�@��\d: b�"O�M���%iJ`�zh���s�'�1O@4��cUv�4���-�*zI$�"O�A �!��PwÀ�L.t��"O�0J�K�	FO�x3�͖0�`� "O(�;�f�	m�����*#��<�'"O2�s�@מ�&����D�!�h�"O�LS��hwh�a�g��] �"Ob��R��4J��b��jp=�F"O��(b�Ü�1V-�V�ݘb"O�����!8-��TㆎJ�i@#"O��`g��PlA��^0ހ��"O$�8�吥_r���r msѪ!	%D��[3�T�.�֡P�`�B��j��$D��`��1t�l����;M��!$D�rw���.�x�狗PS�p:do&4�����i+t3����*�Z��H�<�G�7@������� i,L��4`�n�<�1�V�@����?Q�]u�j�<I���!	d�5o_�/x���qO�|�<�!O8uz,��Ģ�K'���b_�<)�n[v��r�ȞF��8�� w�<�Ĭ�"b"\1�� �p�D�s�Y�<�E/nxє�ۅ�"EQ�*�Q�<�d.��"_��`>t�&�(RaQ�<��+=!)��$�ʑ0� `�c�<��P��=��!R � � 1�Dg�<�W�T���Xq V6+8%v/]�<ї�ۨrE����U��~�cP��a�<��ȓز�ȵ�E) ,���.�[�<ф� %v�JH�k��[�׊AZ�<���$<!�ç_�?�R����U�<���2����*pF(��U�<)�bұp\6�!��'�
�3���P�<�g�C�@XL2�I��]�ҹ��-�t�<�Ꙋq�����+]��%T��y�<q��E�M��Ô��(h�J�AƇ�s�<�+'!8����!.�<J��Gl�<�s�#h�9qf��N_��P�Yp�<���\v��2l�t�b���*�l�<�U�ݹ H1��䈀���sWO�o�<)�"Z�2<z�8s�<^��i+7�Q�<i�m��aM�1�D5!Y��9�MJ�<�@�C�3�n���h�%DwH���eIx�����<�W�MJ�ܪ�%P!A����3��A�<c8V��}�ƅ Z��X)��}�<a��X&/N��wG�gE<	7�y�<Q�/V *`-Sw��M�BBr�<����+p�!
Z�X 
Co�<Y��%�P��m��J˴��$AF�<�dl�jIZ�A�L@�s8М�t��E�<v�6L-�T Ӣm�*Q�І�V�<I���yd�б D�A��xTBU�<q��B�nrb�3� a��K�<�B^?OX(�Fo؊u���^�<i����K�G=pA|�'@�b�<qAf��!�� %�&Y��V�<y5 U,o���2Dlܹ6+����O�< Ĝ�����(:m� 7(Ad�<I0�W"^I���.�X�����c�<����8	yV�B����f����c�<!á�s�4�"Y;`x����_�<�0O�5;�,s���l}�!��a�<� �pQW�W�!g���U��<9!"O�-�DF�.]7v�'16��w"O*@�v�Y�a��}�L�����U"O �@a�ԵC�ּ��,��"M�U�1"O
�c�gG$d��RS,��D/���"OJY��H͝d�jL(P�S1�V0:"O �I�)�$�r͉�B�s¤q�b"O�](���w�xl�C�DN��"Ox���,U�D��)�EI"O�53���>o�U2Aݗ5��I+G"O¡c�v�M�# ޲�d��"O>}[u .��p"��űC���0"O���/:a�l:u�.,v�$�F"O��u�]�i9x�q��	ZS�l��"O�� *Σ66��	�.R�"O�ر�i�+�(`c�M�3�8�"O$ض�Z�%4���'jp��"O���%�~��<J0��V�&"ON�)�kW]��K�KF�{����"O�!�!���{ڶ��J�-w��Й�"O|�)�ֆY�T�Iۧ'{"��G"OZ��#���L§�8}�"��"OpQ1��*`�`�ڔF� 2�F"O����Ƿ~��mń 3X�Á"O���FH�$.����	U�Yld��"OJ,jA�N���K`H΢�hT;G"O�Җ �w��,���_gR-R"O&���\)���R1��+[6pt"O��CwBK2^=�`����2"��#�"O��ᗢ�2��<xŤ� ���"O��[fn�=Z7���dӌ8b"OT� ��^�1)<I ����r��"ON�:�ƊZ?̱룠\�>f<3"OL\[���#UP�Da�n�l�p���"O<��`ɑX�+��0}P&�ڄ�yr�)X*I���Հ���b�����yb�
n���3񀎩
��bT�	'�y�)��;1�981�_/���)�'�y��Na(��uN�B$]���N��yRm��f�B�;��L	A��T���y��9��2�[2Mx���+�$�y���4T�LFbBG��{�����y"�قpp]-��B&&��Ҋ���y₝#6�(K�C� ;�H���E�)�yB�A=��3�&d�������y���2��\1��[����#cQ��y�㞀>��1`�CJ�13����y¤ʯH^P$�V�,���@�E���y"��*�����7&�3�ę�yb�j�j���z�ɂe�P�y"�K�0d���E]hP���ƪ�y�,�4_efU��o��+M��9�L��y��J�&�)XWL�"��=Aؘ�yr)�7vH*7 ȍ(��B'l\)�y򤎄7��8�u�B��P�֮X��y_�~�P�*��l�z����ybHJ�HQ�P���
~���	ʇ�y"NX�	��i�W L���������yǄ!Y2I3c�B0�$̈�Ч�y2E=9�B���}��q��BO3�y��#l��\XT,S&�����#�y�@<&��WJ�0i��$&�&�y�"4w��E�Q.��x$��0�*��	�d��r��<��hK�%@�7z���S�? H9Yp�T*i�h@x�<}JT�%"O�h2!'�x[`t��!�p:�"O��b ��uH�Z4�W}eG"O��5'C�<����v��-�:���"OZ}*�޴>�p��  P���"O�<��g5x@ɫ�ˌ��(M�'"O��#K�J�D1gj\<��E�$"OhIˁgL�
�zxc��+`yV��"O�8�Cͮt+�]1�g'aS�E��"O.�j�e��o~�pЬYhE�@;#"O���)�.l����^y0N1��"O]�T�#/]�p�EA��k"d\�"O��p"��:�&���.��dF�Yu"Oѫ�&ƀhd8����1<����T"Olp!"�ۧU��@yƪP�?�.�Z�"O~a��� ~��������ɤE`"O�PC�b͸(���v��91'r@&"O����1D��<�E@>�@A"O&�R��	���ـG@���Ł"OXq`��ۓF�.%�'�� ]��
�"O�͚�W*KWހ��%(�I�"O��;t
�s
HS��آð�c""O:�;.^8����Nͼ]Ăѐ"O��r`F�<V:��y& ���>=�@"O� S��
�p:�[UO1}�z\��"O6DKXS�9W,Y��(�
��r�<�$+<`б�m\��ֱBF��m�<��ő_8rq¡���Y� ��\T�<�5���!�0��6��y��.T�ؘ$i��k��ȡ���W����A�<D�Xvk[	P�H�`Nْ//$=
6D�p��O,_}��*C�M���r�H1D�� d�|���8�O����j4D� 1�I;��p� )ې���$�3D�"�Y&IX���uN������ւ2D�0�6O1l�^���Eձr#��rWj3D��`��ݬY�.1�R- 5NA�1`�'2D�ٔ��P���Ϙ;���+v.D���f�h"4� �Vh�$83�*D�<������R��=�p�+D�t��Lѽ,N��z�ܾ��A�dl+D��A磁yj�k�ޭ>�-9R-D����n\ر@��?|�Х�8D��k�L�?J�i��[��8á�6D�|Z����j�8�ȣe[fVp�h�`(D�l1�и2 �L���2`$Y#��"D���EC	�)��I����*�q�Ą D�Dq�ރ4�~̩��$tMbN*D�p�&����#�A�d1>IE&D���@X,3���&�B�`�Bb�?D�t��#+�P0$��+�∲�?D���U�ɦH��	�TΜ�3?�dy��<D�p��5|��h��\F��"�'D��'�U%.�9�MW�X�8H+�#D�`�#���p��q�Ӭ�>62LD��!D����l&y�1��EW2�l�A�� D���'�ɚE��A�ՃS3���0�<D�\Ȗ��@HmyuJQrn*@
Q�5D���B�	P�r )�a�65I���2D��#e�v<�&㒶l3��rN,D�����6!��ӑ�)ݰ�@Ћ?D��"�
�Vf8��EP$j���.?D�\�k��YMN8aւ�Ӫ�@�b*D�@�(�*����+��0�^�7�5D�� �y@�
˜\�� �CIY(�����"O��f�]�o�:̛�HO3G�\��R"On�S&�v�� r�%U�M��$"O�p ��E:sbn�[�.Ş1k53"O�%��e�d�5�C�@�H	ĚW"On�"w��`%̙y�Sϰ���"O�5!u��;�� U��.��#"O.P��dG	R�2$Ӊ ��e"O@��b_�7N�'�<GئmKS"O��CE��[Aα#&Mk\��"O��R㌴U�j�)`
I�=\�(��"O�4���9S$`��H�f9��;�"O�U�'G�юH��cW2mB�"O��
�(�!�q���,cDF�"O��F/˭h�JƓB0���"O�4jRJ�-S܀���J3/G��S"O6Q�E�@&Z$n�`f�� `T�S�"O܁bUkҮ2B�9y�d�N�HS"OP�0#iG!�@#�,];{Bx��"O�ʒTd<�DL�D<b���"O�����^M.���c3��k�"O`�ㄦ	7\����7m�!jҍ�U"O��`�P�j�\��KM�Wʈ�"O��C�JJ%]l@k�)� i?Z͐"O�����Z�C7v���A�z�z��@"O�<��C�GG �	��,r��"O�\R�g,�4H#����E�L� "O"���ׄq�P%�@������2"O�hB�ŷF���QE�P����"O��h���	|���p��@�8�\�y�"O�0��I��A(T9G�d��`�"�yb�jvl q��?	j���@���y@(v��q���6~�JV(դ�y��҈K�~� ύN�EI��K�yBnE��rU�gH7u�9˖� �y� }-�袢	\��,�7�O��y∃�"j�8ۓΛ�^wR 'GH�y�)���2���iѣ@�z��%�Ԡ�y2KF�M��	E�1�f����B�y"*U�9r���-� +"�,{��[�y�kԀD�( �h<��3��A��yB���R"��Ӑ~�U!����y�G�ot�Ib�?_޹'�Ц�y��܅Et��B�抖2u����)�(�y������9��'I�EJ�	Ѳ�y�M��D��Qʗc�<#;�41�g+�y�X�6�thA�J��:�B(��yr+�J�����A$E�@)��E��y"4�P�p�v����"�y�o�;l�>�����0�cC��y2ʛ1},��a+�~ �q�q`��yҡ�y�T�nݩmZe��2�y�w�D�QE��hE��.O��y��N嶐����*�H���K��yr�-!A|IQ�V�0��S'J��y"�H�(�� ���=[ܱ_�y�#_{�%�eU88b���b0�yr"�&b3����Ҙ1��LS��y"��f�7I�qXv׫�%S�!�Q�44�M�pOٽ6L�4 p*�r2!�$�*S��IҠ�d2���SDH�I}!��4zZx��ƅ�S���u�$Sc!��
L"@�P�ü��Z��@L!�$�;qO�6�\.A��A�@��!�� ^A��F�/��!7t��肄"O���!�1iq̥�SE׎_.�"O��  ���m#��ƫ'u��I�"ObM8���<I�n�@ğ� i�sR"O�a�#���\,d<`cǗfS���"O�-��!��S�^���!�)0��r"O`�s`N�0LBAI�
��gq|��"O�xB�Ąa���b&oOR���"OΰDǍ��D9w�ɻZH��#"O�p���ZF��l��l�%J�� "O��*+���*5���-��"�"O��bs�d	 $�0��~��K�"O��[���TM��t�˱אݙ�"ORz��9����.
����Ď�y��ڈy�$ppG
(��r�͓��y���[��@Q�$���EM:�y������T�����Bڴ�y)�n��*ѨyxfE��`L��y��\�nq`$��	 `(1ʖ���yb�X"��`�B���81��dP��y��� �� �W��Ȉ���y�g�.!l�Q�`Q�PC�%
��yBd���th�,�9G�B�����y���k���T�?. �"���5�y̐�"*Zd����4e��A�����y�
8q�
ݩ��&)����ف�y�F[�n}���_ ��aq��y�l�"�����-݅�����α�y�MJ�s�v�ҷ��
�+��;�y�d�0-� �Z����` vU
�ɛ�yr��V�~ {UOH�.���ja�@�y� 9,�,���c��9!��*�'�<囤L_�$���9skY+7��
�'���@�nA�3��U"��Ǥ8D� 
�'*���%eաZ�X�SR-�:H����	�'"�[%���f(F�� j�E�p!q	�';�Ea��H�.ܢ�� OJ(;Q�y�'����gaU>@+���gg�����'�0z�d��P�T�ɧ*�N���'�h�����Q�B쓪	��y��%��f��S��E'���dI�<)E�8,^�{p�4f� �jH]�<���=Ĭ ���L(	�& P�KEZ�<9`�ƨ5A����!B!.�Rx�CKU�<y��i�� �Ӡy�Z�SQl{�<auk�a\L���4s|�Q{���\�<)�]-lȹ� ��n��r�n�<!$k�Cvf��gA\�$G� ڰ3T�\r�B�
�(�B�e�E��t�Fh3D��X�!��������'vl�h{ n0D�Xj$�L�p��bA�;��hS�8D� ��-H4S��P��R�ĸ��6D�� D�Ηx���GJH�28��ꢀ5D��0�gۘ�b���0��{B�4D���灖n������'D�-��4D�3��}��#dL�(8���Ӗ3D�\��@Qd�c��F,��8���,D��cӁ�EdX�T ��0i�T�d+)D��k�<'h(ԓ$4f/��Z��9D�L� k.K�p��6%P"z�t���	-D� �-J&㒵�%!&n�~�#��?D�P�˘^Ud��m�O4���>D��:
�F��ځ���C�����)D��`C��i�y����q�T-d�B�)� �*�f�c�zU(�%6+�NI� "O�Ih��7��cs��ĐSB"O<��Iͤ7LP2cǄ��8�k"Oy�g�UZ�Ѣ$��0��a!�"OHЁ㉄j8������P�*OV|K��W�h�3b�)�<�
�'�<����>���q����6}�'�����+Ϣ`�pL��}�T�'���� ډ)O�u�S�;n�Z�`�'R(X$$˂X�>=��`�:j�Di �' ���5�(�5��	.�T��'���!��m�$T��O�'��| �'�Bt�a&��*��õe�	ƺ�	�'hΐ�1B+Z�dB��[,F��}z	�'u�aU˔�gPP�De��,+	�'l�� D*��E-���P��'оm�HX�.�"Ase,"T��	�'q�l���4y�&uj�(��	O||Q�'.��t�ӫ(�E�,����{
�'���8&�@4�BU���H�	�'�����Z%!�aB2�Q(	�'�H]���6Aj��qNʨ0L.P��'h�-+%��=eL�r�K\}�t1��'3�}�p拢6ln�q�k��d2lY�'~�˴�Ě� �{$�ث_�ؽ!�'Hv���mQ��pp�oZ�Rn 0�
�'��Q�.Sp��A���V:�9�
�'���"�N5[V(�`�J��Ys�'$��g͑j�~�I6�$}����'���0B�J�> ��-S	q`h���'lh����Lu����&5�����'ѐ1�g���h$�
Ua�50�o�<�SM�z���(���%_��s�f�<��`Q�s��Hc�N�o��+��_�<�5�K0�yq�
E�(x��b��F�<�#�
2��][!�F"�~�v�
}�<їkL�q���y��ӛp��!��~�<�emL��F��"��,�:�;d��!��/��:�AͲ�B�{�m͊B�!���W;h=s�J�=y:��&c�<}�!�-g����eǕ9�6�1�ᙄ:z!��*_2@P�ǱX��Uوt!���FK� :'fىM��Tul�z�!�d�R�����N�x5�\�Wl�!�$ٌ%] �f&ʐo'����ȋl�!���0D�Ƞ+�+T�_}���b\Yl!�$]<`��#��\�������Q!�$���c��΃]䂵*�G�d$!�d��Y�^0��� :�BD��F@x�!�$W�M� ��Ԓ��t`����!�d��E:��s�#+%�&��-?�!򄁄
������,��5�ģ��!� J�z��Q��8|�JT��4�!�D��V��b�S� ތ��^j!���Zwn��(\$[������K!�!��L�/�����E)oZ��	_$:�!��9tD�lb"@ĶiZ$��*X�!���8Z(�%��.]�:���%	�s�!�D�zRA�s��
�������z�!�dO�8���(ܒ<����$�q�!�DU+*U��-;
&�d�k�lx!�ݴhO���iN$	=��i��� _!�d��8���F�F�Lr��-�!�]2~EܱZp������ܢ*!�� ���E��#4��e�! �d��h(#"O�գ��0`����	�A�z��"OZ@���ц?L���P-��kFb��"O�q�k�=��푰��8*1X	��"O��8�J�cS&��� ɺIu^eX"OnS�˝,u�)�� Yrm�1zt"O(�C�+����e`C�rk`Ei�"OD#��N�jqQ⌋%/ex���"O���1ʊA���3)� a(��"O�@��,�?B�YR��MK���"O������`v��
 ,¸a�"OP�&� {=N��Dڶ[��0u*Oj�K2��&���˦�q�����'����g�-Ɍs���%TQ��c�'�@�bd�k2Ԛ�OԸR{�4��'�h-3D�*;Z�i�憕Gw`��'�&ቢk�.�y���$?��r	�'Op �c7|�^4S�b�#>�>�x�'�y1,�;\t���/::vv0��'�p��!��2U:hC�m�2fNt�
�'"@Bc�z`�U`*,L��'����f*�tM.�*��)��)��'�<Ly0j�-���7%ژa��'�2U��.��oR*aH���;����'�PPk�l"&١����P��'JL�3ƃY����@͇G��e��'���c�KS-*�2%��HJ�*�H�A�'"D2Ѥ���=����$�����'�q{���>D��;piT�N��s
�'z�xŧVx�	�G�Q��Mx�'� �ՠN�/�FD�'&ا����'��3#f�&�U��koP���'��s��0bpY��`d��'���R��~�� 끨����'��W��.
d(��(��d�J
�'w��"�H�ڭ�E������'���WZ�X�(@1Ś�~t�C�'���ɣ���8D����}6 �0�'P\�� mC)�$���E�H���R�'FJE��I�&�@بD��
��r�'y�9��C�9|`���
C����'@��%L@�Sg�J�#X|���':¡����<
0E�#A��#h;�'�F`����t�	�%��^�6*�'������`x�+�~�F}��'��	�i�	���h����x�>���'�dX'ΉU��3C�s�Xmb�'��f,�$u.�	�k@�X��j	�'<֍����B�~Y�գH"R�HP�	�' ��[��'v�+P�O9~��'2(�[�",GY$���9I�q��'#4��b A�/�����ާI���
�'�X��jM�?9 ��a! �(��
�'�b�8U��{f^Eŏ�-H�\��'1��A��@;'y�pu ��T�z�I�' ����?m�T����զ4��%`�')>�aI3E����e/�/(P ��
�'���H�L�-`<��S$kS"�@�
�'v|�w��VQ(��MJu\i	�'J&X����e��)IIѮ$�i�	�'��!��I�?}��G!޶ ְ��'W�`Gh�<zX20a0����$� �'I$����M�f^Zc�� p��'���1�UĐ��Cܽ^�u�f�)��<� �x���3F�,`F��,RE�ib�"O~�U��*-lD��N�`Ԕ�2�Z�LG{��ic���qD�Y{�L՜y!�DܛZ,�1�WC���#2�л#�'x�|�/Y�7$a���F��6���yb��d��l����!J�<�ք�y�ꅒr/�!�ɓ�Hw^dY��
�y��`i(�X��/D�<0a�ދ�yc�L�~@�]%%�\H�H�8��C��џ��Y�)�IZ5�N���,�g�%D��QwS7�N|�wꞘ"����m#D�ԡ��kr�݁�M�&�.��Ѐ%�q̓�H��H�'��*W`P�i@KJ�Ld"Odm�B-�6�r��A�+N~�Y��;O��d��i�O(�B�
l�fr�_�k���(w"Oz�+'�"���E�_6S�r��t�i�ў"~n�(O��qH�C�(g�
�c�bխ)��B�I�K=�YH1ES�l3D�����M[�'�ў�?e�2D*t�x�s(6���:2�.D�P�r)�hvDR"=�,\�A:扖�HO1�z��EC�����G	i~��V"O��P�F/;�\���؏�+a�p�<�	/��]�V�]�$��P�7eOiy�'�
4�=�����x��x�����h$rMąnu!���Ϧm�Q��&�r�Z�
Z�K��@�d-�$�O����::�V�8�b�B�����D\� f�xb剠+��u��Q?BrT���i�v���*b����%E��t�s�ۻ1@�'�5�>����?JS�l�h�8O2ja�`nX�ZY!��և{C�9�T/�a\�aC���+>��'�2�ۓ:�ĉ*mK ����/Z�V����M;�&��.��໦/a{�\���Ax��FxR�"��x�D����1Pt���0<��:0oty!�^�&{8��5�t�C�ɯRI�I�u)��_�,���Ɣ������ORe�{��)^��%���Z3
Ի䡓��"B�77�][�Lհm�4|d*Q#&������7�	s�'�Ľ0�d�a��2��
�%g.��'�Fxs.��=s�e�+�$�XěL<��,��e�g��?�L�[�&F�0}��Z6�j����f����۟0�`)�ȓNm	�͉^nࠋ7خ��<5����p���Q���K�Ob��0=��L�	=��e#6_�	s!�Tq�Ix8� ��O�]�t���~�\���5D�S����҅�Įܩ4�D����4}��w?qH>���DO�Au�"�V�9��=�\��ȓa�bTB�S"kz��Tn�NJ}�=�ۓj������=I�L�{�`�L�>���Iҟ��'�fFU�ٹ��"J`|S�Kޡy��˕{��q�a>aC�e�6gN3D�!�$F�0L:���<bX��V�{"��[=X�-`2��S<� �!G&��B��<�~ұ,=O�<�ç��gs,Y��Oa��hO�O
0eQ�N�Y�4����:S��9�'E�P�Z�6��$$�$?�2��	�'����UhA�HVdj�h@�Ce���'䑃��V�A��{�BM
:Yn3�'2ў�}2RgB�I�5H�ܹ)촙���w�<�U#�;n�>����	3[�H�CJ�q��"�O��GL*;΀� 垵/@x�:�"O�q$!�P�|��fW$#0ճG"O��H]�Z��T�@�d�0<��"OP��"%N�7s<�ɦCԨRӰy�"O� J�q�MW�V�p���ɬS�nx5"Oj�b �H	|̺����K`�<��E"OJ����[�J��t*
�U�����'�ўp)�JC������Ӌ��Y��4D���T�+�bᩂ�Ҁx��I!o'D�[�f�M� ��g�Tm^��r"q�ң=E��4[�X՚�D.h`� ��!#����F-+�%�.P!��LS��'#�~K�-aJ��4��/���1�0�yR� ����	�X!�l+Dn��Ol�=�OZ��fĳQf��gZ�#B�+
�'<��B���zi�8!@jMG��M�
�'1^a��րM����U�>��t����hO?���!��b�8	)�퐛2k؀�w(Ht�<�˺K�v��"Y�$d$9��Y����'�-@dl�wCx��$�[�QQPd
�'V�h��& $ �¡�KBY�'�,$Za)��b؜��(�2G��	�'�:��@$T)x=TaH����F_���7�3�S��?Q�邀b�܈�抙"䤩2��K~�<�DЊ*��9A���"N�Z�j��Tz?�M>��%a���#��q1ԔQA�&R�D��I0|���I.vn��ɱ�	�U�x���'a�LC�Ig<B}Z���lw�0� �/�B�ɰ�Vx�mI�Z6��~�t��ȓ�9�d��N6�1�`&_8 ��S�� B���(A����GS�����M�t��HR\I'���fެx��vb��ɛ8�D� V���/�ȝ��Z�� ԇ�3!�|a�L�8Ep��ȓ��AUG֟J�jIhu���h���$qA�6�~�PX.�zY��l��cpG��P���a���)���ȓZ{�	�C��~���i�+�.n�2���;L��H�P<�d�4��-&̹��>�����P �i�6J])O�����c4�*fD�{��Z$E]6z� ˳"O�h�@\�h��LrԄ��fg��{C�'�Q�`�ң X����+[�a%���!!Oң=94F�,�`�(�CލF$f�-F�<��Ѳ;�p��ʊE��@!��]?y���Ӿ1
p��HW9(���JæL��B�I0;�&�PĂ�4]� ��a.�!2a���M� %�Ş th�ӊ�!dr�X'������jmn�#~������'���:�!��B�>͘����φ)~:�:��	q�">Y�A<�'p{ p*��7q�,Ҡ��'�2E�ȓE0B$�cK47|Q��
�3A`@���q�	�jf���-H���! ��yT�"<9ϓ]sx5��
Z=cɞ\�\��D/D��CJ�,#���U�7;����0D����<�ε�a��L�\�k��/D���ӆG(T�^�C�l��*����]h<���*�09a�j�!�
�SC{(��d�"���� ¼s@Jl�F啄D�az2g2���D<�Y��
p8t̉&)��B�ɊcX�=)&-�v�0�kD ��B�I�~А�Y@)S*�=�4m��V nB䉇 /�$ ��*4��A&$���<Ot��d�"F�����	#�bA�/�yd!�$Ô�=�W�
�\＜�70_!���[b� tB��"�>��GaJCa~�_�l+��ڰ 
X���'G�𙖦&D�\y�Mu�L�0S�F�6I��"�>D�� Ԓ&CT�3��RgBJ07�1�"O�@��)47"Y`�O�X��;�"Oqrŏ
����VD9$N�`""O2�[5)��l���A͞�%��R�"O��K���(3�eas�6`&�$i�"O����dڶB������%����s"Oʼ�p	Y�g�d�aD�C^�)��"Ov%!V���*�|M0]D�Z�"O�qyc��(�� Г��6M����"O�1b�Ońt��cG�jT$�"O�= (�'B����C�� rjB"O�����%E�Yt������"O�`�G����h�u�H�q�F��Q"OJ�r�&I�逡B"<��Ƞ�"O �aF��'^�����hR��"O(���Q7re!��:d��Q"O:�nľ\��`F@=�jq��"O���i͍;�� t��y~� 3e"O�8�@��v�z=* �4}}"��*O��F\�����A+�+kW�D��'V�l�#R)"� �a���fk�eX�'0��*A�/n$����Kd�\)3�'8�%���8�����J�(_z�<��'t�`���^PZ�H ��V �`��'P: )��	y���wJL6#�Pi�'W� �@n70TH��X�\Ĺ��'.��V�;S��`( ��8N]8�+�'[h��vj�+*k��[+K�U
 ���'��DY�k�F;R��m�L
L0+�'@���A��D2�p��!N�/TFD��'2��V�AQ�H
�/«%�]�'��d��M�5{3Yd퍽S�C
�~E�$�:.����,�L2������p!�ȓI�2 [5�PgB�A!�̮%����ȓ;&�`��Q�(��dg��E����kmf<�SM�c�<H@a�	+a�؄ȓd&0D��Aϱ	�"��BCI�@�ȓ���y�+�$8Ľ[�o�/�Xą�'��h!#*8e��8!�^�VYQ��[�
�a�E�4:���$d!,C�	c����E�Zu��D� ^�
	��\��!QJ}JȲ�)B$w�Rt��M���*���W�"\��+-T������;�FL+&���+>&�̄�:eʸisH� 1Ǹ��2)�)�Vx��*��d�ꗼ8�nm��X"�h���E�y�(9��A��a%��d���H9�D6KR�9�p�ɏJ�<	���*x�]� I6��p��/y>|��ӾA�<���B�u���@�
 7�!�d�0<�h,AA(T��uK'�� �!���t�(��(�8j�u@���S!�$@�A"�Y�A��& 6��0��%%!�$�# E�0���ޅz�ҤR��$,!��Ȟb��p���Z�l�P9���#!��ӡl\�u3'���G:*���,Ë<I!�P�	��
�O'�ipӫN&<!�$ /~7нQ� ��;t{��F!�ڨ>�l���-�#�\�����A!�D������Τ|S���W$	�!��*n���,�v0 ��Vc_�!��[�O�䭩t�n�pi�tc͉M�!�Ā� ��K?5��PZ���Fr!��B���p k����u��aH�!�� ���׳8�\2E�оUP��e"OJM��@�9L����C���!"O�$�f��D���	��ܧB��I#"O�I�Ηw:�
��7<@nX��"O���Գs��4(�l�2dE� �w"O`�Qp��^+�� UN�3�\�"O�Q���/�
����� ��c'"O�iqf�L&e��fؼq����"O�]ЀnO �0,Y�ƈ��X��"O�y腍�
2ؐ������"OHAq��|�zu3�7K�>�>h��tނ zD�.]	�\�3醳<�]�ȓUZ�\xaȍ7�^�Hկ/Q�D���Qb�m��oά]���E�����}�ȓ,j�p��κs1e^'wvX�ȓK��$���RNa��%�4to>��ȓ������E,���O
�2:$��hBE���	I� =Ç�:�Vd�ȓ,?��Rl˩x�`t9soI^�A�ȓ\`6$��Ŝ���NI F��D��gI�ai!i޺_�,ݐ��OX��H�ȓ!?ԕ!�iZ-:z���h�B�M�ȓq�5���#�20�H=L�]��S:L`��Ӛ5
���m#i�.e�ȓ:0V̘!ME�$c�d�Bhܡs����c8����5�\ٱkǙnN��ȓ`���B �^���S� ˓1�ځ�ȓ/8�[fC�Ch�Ó�\�k�*|��%��R`�G7z����	(Bi��ofrI�㊥kZ�#�#��G[��ȓ8�I��o0�X� CB�?t�ȓQ����Ǥ��*�� Xh��=��{h���RA!8�EҔj.6�.���4���H��>���kN./l���:�5����q(��+Ԅ�l�X �ȓco�ܠ��ȋ@�4�s'�0:��H�'F\ "�ɝX���q@/H#L�	-G�jW�����5�OP]���W���0�U�
�b�����p��%z�Pq0��-!qO?���"�KW#Q�\�����>�Ov0Q3Ώ�0c��S lĘOe���U�+Zc�B3�	~�b�8���^��V+L�[mL%���'�h��7��=�����!̤9�V�x���s�Q�.�����u��^hl��cD�ˣ�ZX �&���5�JI&�.���%G�.����*M;�y"K���*Yq��+%���ۧΚ(;���,�$%>�:b���~��+@��$A2*&������~��>p�u��5)�3���F���*�`ʛ��9�fmB7Cd�Bm�1 ����!��,��暐-�:%s�IX:���a xn��b-R1�����}�$I�Hl���\�x ������'z�fk�)C��� $V!*������m�������p�H��l*Q�a�(
���L�QC��H" ����%A�5�"���ϓ�;f ����	K͖�
nÈ,�2��#���\[H����,3�8����9r�%��eH��v�0�%D(y��u@��pl�0Q	�v�',��ӶD��	v����~ 3aB-.�0Q#4�M�`l�o�b$L ��%%h���ӌ�y(�Ƃ�_VѨa%��X��q��R�XjsO4�	)Ƙ'Ċ�����+C������/�������Y �r@� �5
?
W�Dɕ�ߨ�]i OP y�
� ŋ�_,��J�a���I�lt�`Ò��+��`�b�+�,��V���ٔ�?S*�m�cMO�iR�ô�VIqH�#u"_�>��d�T�Ϙ�N��Ҿ'�4�FJY�ɕFD�Q�J�����O��ZF�'�QjSh߲J��@�QK�n�;�ا0������wT�٤�G8f�M:�Ȟ1L���x��ќJ�b��wM��9�
J�<<�)��R�v}{�$�S�arJUt���(�
2}�n`���� M�B�9���t��8�7��ƦmX 	V�>�d���NSb����0Շ�~2��[�Nɣ�AB9;������ܜeVQ��Qv��>� �h;�R;<��p8+_�
�D��sO�(;�`�s3�>Or��P�T�9�����ֻ4�@��4��8����~�1O�)�u��Asй�p*͜7�,��лi���O��Y�B�����Bvح� ��5�$����ܳ[�Mٷ�wqt)9R)Ϛ5(	@�����5j���`��9�!��Pd�0�V	�-ВY1V.˟gB�8��#iw����Y�`��)�a�Qf��S�?J.Ry���SlO]Z�\{�%]�K�">�����DE<���%hF�B�ˋ>C7\�SDbj`9i��*v���oڋq��|
M�'L��|� �\�wI�=�t� ��S�^J.����'��"=�O>����	����2I%=�){Td�0�Xe���59F���S�ѲF@:�8�K��S��F@��7L �z���Mk�����Kw:ʓ .���?:��d�� 	�X,�c>q���\��|��.�f ��)�M�/9,�'ڒ��4I��Dy���h�GW H �m�F��)X�0�Eކ9sr	�4�^�h���?�&?i0t�?}���ӧ[	8G�����ě_E�l8� ��=a{�(�D؁P� �2���2L��k3@Y�(��əe���h�T��;`����0���>�'邕�s�ۄ@�h!DDQk����hO�>Q�ׄ�
���ҭǀ.N��1 j�OLő��
-�t��D�<��p%���� V잌�é�/ߒ�jY���]�����(O����I^����%�p9��O?�*	M���EȆ�=sў���'m4,���4?1<�Wǔ�X(x�'aLGyJ~b�%6j:4��G��b��jv(E4mX�����~f">9��	Q�?/ �/ĜA��L�7>��x$!Q�y��>��%e��У���l>�S��S -������ev�{!@����7��|ʉ{�ǂp�څ�g��/!I��S�ʍ��~�n�<_xO.�O]|�|"c��
N���q��4����M�H��hO�]�Ȣv��!d�R�r�jʿ@N������O�7��]�R��Vy*��OБ9T�
\.�0�#,�ԑ�!�IY�'<�锡d�t��e�8fN�u����V�����?yr�3�X���'~�ĠV�;al5bЈ�?�.h��',��$?���'��mŉJ��Xy�cЫrU����:�yrA�:�Hqd��s�4�ʂ�L���h�nԕ'`����|�O�S��ʭ��gI�12�٨1�˹KԼ���Ru?A�m\=�����˪Ю�+Q�̦���������ƣǉN8L�΄����v�XĨOx�lZ	C��?�xD��
$z���ſv�4=�rl1�����5���:�Ӏ�,��؂@���h���\$�d%��?��	�Z�����J٨f6z��tN�Xq"OP��5)�P�ؔ0OQ�N�ZI�U�>!q�5ړ�U�aW�p&VH0ê|\�ೳ�'���2Y�Jc�n#~�������h��hO>�� �P���[�"�kƼ��2��ȟU����8T5Ҁ� �@����"|O�i9�ā!3�IQ� ���2ɵ�O�=E���		R*<�L��D=��Q�NS��yr�ڱHbTy$�Ԅu��	XS)Y���	iX�({��Q��@�bΚ-�pj&3���O���)�t��`�S�ܑ�C�3w�b���)H�!)_6���M/@�����7Op�a� ��:b��R@lˏ]�$kCcUO��������bZ|b��Ɨ9O���� g���,9Hc��tŎB�I�P��=�Q��[gLa�r�M����̘�H>qT�L�J�"A���X5L�.���' Z-��*�P~�?�&>ip5��J�a#b�^�b�~L���:?�.O$�O������@T�x+��st��ss��Bd�F˓p"H�4L��	(�'>c��J�震@%��"!LS!TÒi���nyB�Q'�M#I>AF�M����C��&}���S��U�q�0�X�>�>h��M�1O6O�ʓ32��QÀ��=�68�� X�'5�˓�~2#X7
x���o"B���?��r�	�oV:��A�#F��B�-}r�x���).є�k�E��A��XI$g	5!f�;VZ��!4*��BxȄ@B���S����O���Wh� p����3$~���f�Ĺ<�������'�N�Z1LՓW�]n�m���������'�t���J�N옖_>�c�2* �O���;n��y�W�ɖ�?��@�.-��N<����-�L�3i�1k~�i�D牶�(*��W!�(��f}R�'%�*Ï?NEHlᦩ��b>b츮O�y
�K6OW��5�M;Q�=JKVX�^�~r�'%t�r!�c�`Pq��D0����&�'�8 3��[-^�XL���y��`����8v�p��Bҟ��IM�v\�GImN���4D؋cO)cZhm(W�\�.�NaGybn�70P��ώi�OV��'��;�5K�eK�j|���`�N��K�|��hy�- �f��P �Ңv��!`d�VRn�a��^  <6:�n�^��?��J|����*���BasP���Y�bd�D��/�H)�#N����v�Eq�Mj3��x�5·4$#֐SW�>��K���[O�Tq�͉�6��p�F�'��m`��)�O�0�D1!_�� fĠsl��Q�^u��b�D�8�cC�Dѝ�M���ԟ�ɰF����q������A�0�6���,��$�2a>uXvȒ7];����&�[�*�"�
U�I�%�p�i�&�8���Or�a�Sut�
Q	F�V9!t J- �˗):8�J�H��`�������ē��D�q�R�>�����B�	�Z�[G�-�ORXc�N���	��B+Ue�� EB�9E�Y�T�I`;.�ZE�^�	U.�C�O��	�ܠ� R*"F��)؃0\H����&`�x1a f�(5h�ց8F`��Oʂw���X""O@��嗰k����ZMݨ�A�	���?=ɵ��=$sb���]	E�����i!ʓ}�����V?DM��އa  �k��/2�����h��ȟ�ػw���yb2aX�@��٦��=�Px�k�/����*�36���1�j6�� ��ɨ3�\$q��G,;�`@����7����d��~��KV�v�`#G)�h��b ��yb�#&�Q���s�H��'���Of���	@KXbaڱ���Q��)Vl��@h!�D$@��DQ$	:��!�K��4j�Ɍ$A�S�����S�OBUY��G�]f�`��p
�'��誃M���f�p��)X-��
�'�����E]�����IF6Ui�l3�'%hr�a���t���8SHV4q
�'� i�!NZ>�ڠ2��� Bо�	�'�t���A�[h|���_Jjqk	�'���B@ԳC�Nԛ��03��x��'�"KҬ��N������/5����' 6@p�鑹�dQ��ʈm�hj�'tZ��2���.�ҭ4	?�%z�'A�h�I�	��(5�F$hl��'6��ȵ�_��H�05-��w�V���'t�0�A�&$D᠁�B:e�0��'��؁�牭9�>AaQJe��͂�'!ڠ�A��*��{VCD3`�"\��'T��8�XP��Y�6@4t��}Q�'��]�D%�pK�Q�����h2�b�'R|ī�'`������t���
�'u(�!�:&���tl� fm�	�'��	��]:�*P
�M�}ڂ���'�����	���bάa��U�'@�� 村,P�	A��1Y,D]�
�'����
�z��x�_(,�:�+
�'xD A��K�J�D �VSR�	�';^�Cs�ٙ�H,����L��H�	�'�3E�J�)�N�)�_q�2�y	�'B���|���ڔ`�tx	�'��h{�F�?��*AB�o(��S�'�>��F Q�g��Сφo����'W6��ꈉ��a�M\�cy��(	�'��("�
ʹ�����]_0��e��<H�H���L}��#�aX���~����2��0Yt�B��	 `h�ȓ&��)�1�FA#mH
[nJ��2EV��e	ݕ- ]�E��<^�T��e����D�l)�`��U9x�ȓ2�r�SҦ��A����c�R���E��G=	����
[(������ݢM��v�bە&#8`d\c��$h���ȓiS�� k�^��j1�
趬��EMB��R��?d$Y�7o�%e���ȓRj�DD�RJ�4T�`$ۉ!�~Їȓ.���:g�L�(��8"D�^Č�ȓ.K�Pj�*�,6��i���9{ x���ZZ����И*��x�*S�9
��L��A�!�-9Ed)���ձc�����S�? �D�AꔏN~lІ�ƦH��i`G"Oܩ�e޽X��;��73����"Ovxa6n[k<!�v,��1.����"O�)�	ڵ'�Z�k���x8q�c"O�d@!�V$�DW*n~����"O
U�E�,5�-K&�(e��!"OJ8����-��X�&��"uPR�"O��Ui
,	<�kE��M�Xɦ"O`X0R@ց)�dT�#FU�?"�H��"O��×1P���`Th^�r0t�S"O@�3�K���pv�JH}j��"O�=	 a�#$Tά���و�8�K�"Oz��3Ξ�Ŭ����U1h���"O�H`��S��E���v���E"O�D�5��S�}˥ȗ�U�>	�"OvK�H/�v��׼9�	Qb"OD�P�ˣL4�k��3�����"O��pA#X�.���Ԫ��n��H3D"OT�(0aͰ;�n�ɗ�f<�{�"OH(�&��C:�aɈ&nT	ۓ"O(�#�*O�n+^�������"6"O H� L�NS$�Xb)��d5pA�4"Ofh0�&y�<�R�G�a28�P�"OJ5H�	������F[-��Y�q"O���sLS�hYj�JW��Ūd"O8��#iJ�E�ڡ��I�("B"O�p�R���2f�0z�p�s"O���AdB��T � Q�4"O5@�T�(�(�9����t��"OT�@��2
�c2N�%u�� "O�還 ט{L���:�@q�"O@2���R�`��z��H;"O�y�M�
i*���Dx�a�D"O��E�@�S��
��"�fDÓ"O��E��}���q�i�9�"Ј�"OVT��Ɠ�|4x|;V)�>zp$��"O�l���>'R��7"[�:n��Q"Oҕ��&�2�ЃhƼyTV BD"O�}X毉�SJpĨ�G�J0J`��"O���a%$�!@D�G*�;"OL�C6C�V�b�Pw.y��4��"OK�,�&QH&�\�oy��c��31��r*�丧��R@ɐ��E��Γ�Z��9���y/�4#�6m����M�6��r�Ԭ�y�)ӷ*�и�d�'M"I�P�0�ZP�3扐h��؈�dR�S��)�4;a��&m�O ��Mj�1E�T�_/���1�Ԏz��C�	%���$�����6��;NB��	�'��a�d��I��iR�����MG�� ۡn?&���N�&�0pS�G���x�����N�;6�� E+<�Kvf�!M�81�#)m^؀B�ӹebh4����:4�b���W��>SA�}���J��9,O�u"�"�>�`��� �1V��<���'3��[F[�wy� �Dᝪ	�by�AÛ;m��S��'Qڝ����j*�x7#�6'��P1K�PP���nI`��
:Ȫ 20���l؉&D�/a����m�q'P�V�8;3��dG���6&ѧf=Y7D��j�;ʚ�P�#�ylX���U,*����c�Y<6�V>�z���c3�Һ,q\�*��T+O��D�sJ�3=��$;�h�wD7g�1�T���7�\4�0�G�uJY;6�"J	��L�1�p�b��4a�c��B�.����ad��k9!�j;OJ�F�W���$(��h�Ή둤�0c�2�p�
!W*@h���O fFB$n�<Ҥ b��'zH	 Ɉ7)� ���f�L�i��2o��c䨁�*xy1�8P���]3A���P�r���A2��;z�!S��u!�قA�бIP&)jXh#�U�H�
��m:`LHp��z_q�0�����>I��_4�iZ��4�N�P �VQ(<�P�F�Z/��z��fL�U���N O�%��"�.t��I�����$���O�����z��e���_-bXd(��'�$��"�C>XΠ�p�]��� �����\3P�r���/�nQ
� ��[�J�����
:QP�ڨF�(�����&��'� ����'���+0E�0+C��z�ݟV�D�(�d̩1�-��(0qeH�R Xt��'�0�3�
KqՖ�O�1���d�{#\u��:��'/k8DP��1s�<���̗n3�C�6>�`���J±C�J�yP㊫f,�$�H�* TD��)�'5�#�Ӌ{�h�iA`��/�MB�'��mR�g�n喴���.��i-O��kR�-�X,Z�	��0#���K�h�+��3e<�����b(��`Ȳ��CsF�M. i�b�]�Nѣ�OT�Ћ�w:�Z�
�qR���퉻�(�Z���L����E27J�P��������+�����"O��0�חjd����wiD����'mpa���x�v��O?��4 ΪXT���7gC�tfJLK�<��,��	4��21X5a�k�Ay�P�{��H �nX�HP�ʓ�����[���k��h��}���k�*4P�I[�%���m+y��0O^�`���ēR����jU4D����fm�PG|B�4;e��0E�	G��PUs$�)jZn13�h�:b�!��@���z�Z�{�,=0s�\&'@�DW;!�Ի�{��I��r�2��&�2Ɗ�I���2rJ!�D� ��1m�F����l�Y�!��L=V2Й��ɉ���Dۡ�\�a�!�7n>���I^0[����ȋ�Vq!��_�$z�1#@Zh�r[���'�!��[4ɮ�:T���*;dȡ1G�#oe!�#J��'"ӥ����H"UD!�d�#`��bd�
1Xp	3�@TGF!�
�=1D��F-��z7��
���2�!��7N�V���|;ؕF��;E�!��4����SKI>���C��a�!���[��K1Ǝ�!/�%���
xM!�@���i��T8m�Cw���@�!�$X�@��P`�CH�i2Ck��w!�=A�qd�K�k�X�W`!�$C'��ukU���;�HcU��e!�d� o����%���;�̡a�'>ĕ�Q�W�J��#lRNP�)#�'��e�cnJn͠�p��U��X0��'���&��/⾘À���3�����P��*�R49�4	�&ђ`��7a&$A�/�CB8{UL�3Q���]OZ�i6��:}@�z�G�b�,�ȓo�J9P�)�Rqd�J���y��$��<��H@��_�^��4[�� |�ȓ]b������
]��J�JN�z&F(�ȓJꈘ�$��O��$I��޶gZ����m����a&	=)Uf���h-7��$�O��!�Q�ڸ��OP�<C��ب[n��9�@�Rm��'�r	����,`�$�G@Je~tYC�|R J�gtdI���y!V6.x,1 S��Yi:� ��U���?�!�ַ->��h�m(Vݴ,z�ț�E�,x
���d���d�2̈� �M�%�X�'&�t џ8��3c�p@���	ռN$C�.FU2aQ��9�y�MU�`b�%�R,�?L��a�M���
0/�(��d�7��)�'T�u����k�h!�m��P�
9�ȓ&(P����&S�`\�@A �&�B��>����F!�e�M~�=i���1���Ҳe�n��5	����p���O�qO>�B�A��l�d�54�z��#Ǯk� $!p�׾K�a2)H5�����!_�Z����Ώ��$Яm����6?A�`\�Zц)�]�� 6��7Ȁ��8�V�g�����[ ��*F�����$^�v�a��J6$�p��Z�tHFD�(ޜ��і>E�T���v�z�c�L� IP5.� �(O����	�s�v�s���2JS(���	2���ȑ����O��;@hќ�1�1O� ��e�>;����`iA�G��3��Y IV��ӣ�I���S�O*M���4h$2�y��Ik�$ՙ�"~;XI��|��b�I2�qIUO�S����Mv���(}�����T�D�wi�RiJ�����Ck�|��w���t�U4.v`u+ʮGMNq1��^6D��<���@�P�~88�G�UV��yGy��68�� � E�j�On��� �!�9�&������'�t�Zs�27DH�d ]�>�(�lG/7Q�1K#$�0��)��L��n�Y*����S]�H�S(-D�$�󍂵�
�����23֬<���>1v���?b���דk^���jߒKn4�$eD�LT��	�MP頶i|U�k��*=��jU��G}lDB�'���I�+ލp�`�ʡ��o�z(��'���c��+_V�
ۀX)�P�'��@ �JK�����.d�� �'�]���ժ m�Z�؎�����'�Ŕ`�ҚU��jf'*�,�	�'+����*�/��]K�HFr3��;	�'��]�ak�7%����d'G9u
*���'�����˞K3����ۨ}�x�'Ujy�M�|!��@��7|g��9�'���zaN��bŹ���wf����'Cꐯ�7<��p���\x��M��'u*l�' K,;d�?�D@[�'���c��X��s��)`�I1�'�.�� +��C�=q-6��'D���# ��)�s��`�H��'�����T�E�H��,Y�f.t�'0�Ԋpȃ+��5�#�O��`{�'��0�Tu����2�ɇu����'m��e��nq0 �!�K=0C |y�'G�1��k�8���`�U�+�J��'JଳK1����G��|���'�r��4'%,���w,(��e`�'�P}sG"L,$A��*Gϓ&/mZ5@�'�l����#G~>`��bְ$ô��'PLi!�l&UVR|���.~,#
�'"x�rWB�w�8u`��)%v��	�'&�!ao��M��
�D�)}*�b	�'9���#o�`"�z��U�J��A�p��/�L�J�ZpH�!y��|�S�"F��T�ȓU�����3|DJ����pF���ȓn@l}��$'BpyE��aK����,����V�=���!�_
0��ȓj�(x*��͞�0x�fכ|��|����#�O@�ZN�2�H�=��	�ȓ��� BM,{7��)@E �lה]�Ɠ~�rP�3D
(^�D����0�4��G%;B����O�Q>�(�.Tv�i��jʼ`;�@{���b�@a�'�t$��@q>1��"c-r���C� ����'Wc~��ǒh��%n>� '"j���䈀B3�����@���O� $�9`;R�S�Op]8 �z[4���@��th��'C�E�SC
L?�C[�|n:ҧp��82���M9le�7)����l��G�v��'��	�S�Oo��#,��suA�)
���9�剅9���I>��ī�9k��T�A�V�H*Ba�>Q3��>)2�H��0|����M�^͓QMO<'B����]ß�ѬO�=Ҍ&�)�8{����G��<IĹA��H����b ����T�d����/��f�RHI�a q����y��c������ P>��!�	�G�<�[��F�K��� �HN������W7�ɣ�0|�-ܠ#�����1<��Ĭ�`?�%�L?�/S3��)ҧ
�b�9��fd]q1��,=�o,1��d��"����3O�?�[&A�W���I�V+�5��EZ~?�v��O��Γ.ӱ�T�c.��T���u(�����+/�|�Ȕ�i~��;�.��P]Br�O�3�i�mQP��Q����#.��(��M�"�-O��b��S��0|� j��a&�&x,��ك`	A�d����ky�FO%y��/�F>EC ͇!�t����L�% �BF�>D��z�L�(@��%)Pn�4
Tɘ�B;D�Ԩ��n�z`c�%ߎ'��!R�'�f�cQ�ݨ*9*u[W%�.�����'����ơS�� �ǂ�UVJ��'O�a;1'	�<�$�4�7~�9X	�'tXt�a[�q_�۰&,/��h��'��A!���IrD��%N�.$!f �'/�` Cj9��������2ȓ
�'���@E�eU��{�/���2
�'8I��.�
9�,F�R��B�U��yңB�Bq��0u>5Zt�;�]�y�D��Q�bX5�9d��y�a
��y��*o��T��"\4 �,I����y�f$(�j	S�F)/����S�ڽ�y��Dfr�6P�(е�Q!��y)(u���*	�t��a/�9�y������U����5?�b`r)��y� ]�z�&؛FÙ4)nPs��@��yb�Z'ED I�/�)JQS��ŷ�y�]'�A����
}����N�-�y�V�*`Nx{�!w�D�s�i�	�y��z� <:0l�p9��a���yҭ�;3z}�v�`Dh@�TL���y���K�$(�0�@8R���ֵ�y��1`�正�O�)N΀-��a��yr�?0����7D��B��y��˻y}D�����&����y���+Hp����y?���q�Y��y2���oƶ��mC0E\R��p)	��y�dA�?|�=Q2�\�> I
�2�yR'[�ZVH�?�jQ+ï#�y�Ǉh|.M2���@�Z�a2��0�ybNɦIr���41�����2�y��V2]P��ѮN�1�4[���	�y"��/h.����,`G��(#�S!�y��.u����<H%�P�ŉ��y��HN�;5,G7G���$�(�y")4)�1���/A��	X�ș��y�e�o��QZ�h�t�w@��yb�O�Y�xAY��ԛak$��fC�-�y���(*��0X�,]�j$�� L��yr�FT��б��P4U7@�2�y���8���B��}�&�J��y��Ɛ3� ��a�/~J�f���y��/d�8�V�Q$*.�2�k��yRE ~���Eß�8��
Һ�y�o�L���K���n1;��Œ�y�+�9_Z�a�-v�h���n@��y���2El��瀌(����[��yҡ�Sh|$6�Y#�nX���y�a?Q�=�v���H��I�L�/�y�C�ވ�Z��¾(��H)�[>�y��+�4����x�<����X?�y���?L*�I'��, ��qٱC&�y�I��w>��R���H:s�)��y��1%�q9ɗx	RP�g���y2 ;4�����MԮ:�c$ ���y"H<\n:��D�}��0��A���yB��M*e�D@�d�
̰�
Z��y���s{d��YE�xI��L�yr��:���vJA?h@&����y��ȄjAj�&�X�.��Ih�ǔ�y
� �X"��PqX`Br曻p5��+R"O��3����aZ��ҭ}8j�[�"ON�"�HR�v�N�S#�2��Ye"O0���&�3G����aO3>(�a��"O����"��y���Ӊ��Se"Oz�bB�֎MB���`�8M���"O�V�4帩9��\甴��"O>!���F�3˚�0��:�
-��"O<s �X�m��LIRaA�Om�]�"O�P�&A��"�L�b���2��!("O�Ë�P��mb��D�%�,�k�"O֌���9�$곃B�sŦE��"ON@P���� Q�0�����"OR`�D*ރp� a:6b�0��1r"O���#čg��32#�D<��"OR��	'8�xh:���P��|I�"O�,�b W�	��ԁ�;�H��"O�m�fdI>*X,�� �{�"$b�"O�M��+�)��l�3��4[�B"OZ�{'�\�T�s��������`"Oԅ��)��Kr���lƊ��m�g"OvX��)	�~�z`���5w����"O��
�Ƌ�fǜ����(2�$)`"Or��`a+O������J��6���"O�d�&L�q�р�D�"2���"O��B�ٜ.��c��oQ�xQ&"O����cU#ž�E��?/��C"O��A�)D'"��gb[��<��"O~��t�
k�YP��L|2պ�"O~��@#�=���ǠM���f"O��� j�c�TA!��FuK���2"O^��4��"���˂�K�]�H��r"O���@�Ϯ ��(����1?!^���"O5�����8,j���<F�I(s"OT�kC�D����S��<Y�"Od,��]'Ra���O$4 	qU"O�u�̄,���B��N7a-P'"O"�sԠ�&g�űr!*����"O������7��� �M��m'���"O`��QX�X8z0L¤#�XW"O@�q`���V�� �+��He��V"O`�d���9���J�zax̩ "O��R�M&8�鲂
LC �Q'"O��a�L�Y(����y>,�%"O�e �!Ar�V�'�T�d
NX��"Orrw���,�ԀcA+f�vX�Q"O.E
W���(s�� �Y�j�x�"O����e�B�Zu�|���� "Ol�H �K�ma��R��?��P�"O����#�8$��QI$gZ�7��g"O����H�<۔5Qp�S�$����"O �&^�(�d������M��"O�D����=����/��=�Q"Ona�̏�:lԻ�^�Yk�%:�"O��!ψi�eP� �!p�xt�"Otc �ܬDȈ���Y�1�(	1"Ox[� �4θ��2/2�m�2"O�ic���-c.�`!v��5 x���"O���=+��'j���Q��"O4UXRd��+��H�Ȓ�J|�rU"Ob�0ubK-ML^$�'b�X<uҒ"O�6h@6OJ�r�٨vhZ�a�"OP��W��<+sFl�A��
,`�0"O���࢑H֦�V'qb�2�"O�  m+R#�0>&���t\`���s0"O�9�5��	|"<�,^3�^��"O*q��Z�f*�U�b�p�FLB�"O��)EA�0u���.Z;Y����"O� W�_�Kڑ
 �YE�M��"OB����
^�}c̅� =^!Iq"O��J^"Ӧ�3�ʎ�,ȸ{R"O��ɵ��-mV�����L�M�"O�1�k�SAlq�Vȑ/JU:�i�"OV�r��By�C��_�gNDL�"O��b3
Q�CBO(;؂���"O�m1䇸I?.������'�*}Ò"OvE.u�|m���\ ����T�H��y��K*2�[��~ꮅ��� �y���q�`�A��sFHrW�F#�yb(#!��ED���|� �(
;�yr��Q-��
Ǝв�ʬhSh�=�y"���'Ͼ	16K z�> YT
F��y��X�(C<m#F�0&�,T���yR�	�T���/��!\�yQ�Κ�y�뗘������	��B�+�y��-�ȩ{�c,6��(�H�y­�c2<a���>0�ȩ�1���yb��F�v$�A	�-c�Q��F�y�ɝ:�TQQnY:+���#�	�yr蚰	���( ��/���
F��yҫ�� ( �"�����a�%���yjZ�D��k��{]��˜�y"��<(�Ay��^��p-��dP�y�$^�n��BC��V�kf�A.�y"��ʖh�D�	n��Y��yR�ӇKި
(S�:��a�/�y"���t�
DĜ(#l\|I��׉�y�M�)v�\:���%����G��]���-��gѣ!�(mxE'YfP�ȓul�
a�  X
0���@�A�D�ȓ
7P��ЂG�e��e��j�\���ȓ/G~0rc%]��H��˝$N�.܅ȓI����^0@tݨQ�F\x���-��ȓH� �(��Ċ�x�ұ��[�tr��2u���$\��� �Ųv�ߕ4�͹4�m�N��ȓ7��Q�aÁIi�Yq�hQ1�f��W^�� �Ü�%�L9Qp��}\���ȓT��	����[��V�@�a�RX��{�<�@Ζv�$�+�m���Y 2����-)fŗ�& p���-C���Q�G��=��*Md�ȇ�}yd̒�ߺmê�P^�V+!��n]$�g"�!J�"��0���L��D�� k���g�%}����b�E�`���H�HaX�����|iRH�#[���ȓ}�zu[�F�s>���K!~�h��L �p���%�\I����2^�4��)tS��=�`b4�D�&i��p���A�&S�C��T�h�KG,�ȓ?���?F�`�x��P�uV��p|d0	�M�*Uz�h� X��L�B�rb�%�t�p���l-�e��c�.�[��7SP�]��eE�7�P�ȓ_9d�B�l78FQ��bZ<%Y8��ȓ�dX3rK@]k~�@t�7�*��ȓ,
��[�S�H��3L��nQ�(�ȓro������}e��(�`פ*
(���S�? �����  ����$����"O�|j�A	@�F��c��vz:�8�"O|)�4��	[��
7aJ�wj��Qd"O�jǧL"J�V��R�� �1�U"O�ť�/�p �pcY��0�Bg"O@M9b   ��     G  �  9   .  #<  J  �W  �e  �s  N�  ͎  ��  ��  Ӵ  ڿ  p�  ��  ��  �  _�  ��  ��  +�  q�  � < � �  n" �( M/ �5 �; �B �I P �Y �a �g Pp �w m~ �� � ��  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf"O�Ya��=!l���Ɔ�b�V��!"O�!)��Y�fx���eE\z0	J�"O>��pg�0Z�2=�C�A�Hy�"Ob\B��;h�`��Ɇ*���S"O�h�T�ÕZ(jܫ� ��+�Ƚa""O�A���I�{"��qReM.v�\�J"O�I��cR�G�Fm+De����(�"Ov�M�{�Ҵ�U���F�T��"O� ��M�g��l�a��8{�Y*7"O�Z��іh��8`�tm�`�"O&ESS��M�,ɠ��b��b$"O,y0GD�!�<�Y#dYF��c"OV�Wc�6�:�3�	�C��:�"O�`y!�������3-�<�"O��!S��3C����ǇZ��\�C"O�V��vA����EE�@�J�yT"OtXa�Ǫ|�t�2&�ۥF<��BC"O�i�w��&dUj��+,1�4�"O���I�tͰ5���߷O�y9p"O��&�(w�̕Z���
P�C�"O1@ŏΞ
f�}KT��}�P�&"O@%����-Zw*�`C�#���"O01#�m�{�0Rda�#�"O� �	�e���Z� TX�؉B'"Ot�[��*Y�~����4[�h�1P"O��@�K�4Xպs-َbF�ģ"O�-��H�l붼�t,�0F(���!"O�����G>�`R+�0Zy�6"O�eXu럋>���i��wf�%�Q"O����d"�9c*��h>�`;�"O.T���T�`~fM����q)X�h�"O,�YD�#H��k\��t��"O�ɢ%b��/�P5P!m��hb5�%"O���0�φO�Z��k͡1���k�"O�``I�4g$�1шىK�yR�"O6|�D(
46�jf��\��A8�"O�ukg��<Pz�Aa`�#�h��"O@PQ%ƃ^R��p� �p���"O�xjd�j���a�ݾ
L�t�V"O�(Z�[�3p�����CE���r"O.��E�	Sn���
W)^?n��D"O����)�e=!쎷E+���"O����!,\�| �-Z�6xtb�"O ��.X������.��K
�!	�"O���*� �|�S��N ��irU"Ofl0��h=��@�D 5K��� �"O�<kqO�D�
�AۣFj�@2�"O�2���w��"��QL�.a��"ORp�2H��X��a�Ԇ	���A"O�u3o�A�dr�R3�Vy�!"Oؔ�sO]�:��@��z���U"O4�k�a].����E�j	�p"O�1`�	
 ��x1�F�C���XP"O�𪰇O�<�D�8��$m�p��"O����Ȃ0z�L	���K�(��	ˆ"O0���<�*��4bڥ�V<(�"O�m��OE SX�7$�f�31"O�x��R�8�k�]8�U��"O���/�4Q����TdN�lЌ�Qc"Ov���j�3����cč�Dm��"O��ۗ@^�?1�H��ի:�晀0"O8��M�T#Z�h����B0p�r�"OR|q5��*?��ATn�(Ta+�"O��zc��n��w-ݏ���v"O|��u�&�j���?$��q"O~4���7,��)q�V3h���s"OJ�r3M�i�[��V�ZY�u��"Oҍ�dD 0��ER�<hbv�A%"Ohx�  >,jȁ��"){�M{�"O�(�b�Aq�tQR����]���
�')\5fŋQk���M�r���b�'�~-2�+��'4���Ůe9����'��1gOJ)'}.��a��^�F�'W�1�( a��IJ�s�ź�'"D8"�J�,�^P�"�ب@	�'�ʀ�F�9Q�  �����X��'�p�Z�-3�����5{?���'���-c9@yq�U�i���s�'�5��A�g*f�)A��$u���*�'В}�%�G(}b`�e!Эe���Q�'�Xi���2���@�T�^x�a
�'�^dk�D��h�J�Q��B�d�H��	�'o���� ̗Q�l��@R�]� ���'ƶ�3�ʑ�����F`[�J���'��� !L�,Dl�F��6}� ���'�8#R�F!*(@��5CA	z�����'Ϙ�q� ]�h�P�g�fMT���� �ኃ)4�J&ךF�0�x�"O�\��]-|�9���G��0��"OTE�2cQ~B(�b��)��"OD)@p�1�uKЧ{�a� "O؈+1��6$\�s
�<4�d5h��'��I����I���˟��	���ɮv��U�d�H2�4yQV���Y������P�Iџ|�I��<���� �	ğ��	1A�p��	����kL�2�
�������IΟ��������Ο���ٟ��I;1�.��K
+b�`� ����QVD��ʟ��	̟l�	��������	ş4�I�E��z1c&
ed�01�Ř{�D��I��Iџ����� ���� �Iڟ��ɰ_��չ`H���z���Q*����ڟ��Ꞔ������	���˟��	KwD RdL�5xv�@�2��KJ���ퟬ���d�	����	�����ş��I�2��`���!/'�Y�!�GA:\�Iʟh��ןH�	ğ��I�L�Iǟt��	G�<�c�Z33�I
4ꉲ�d��ǟ��Iڟ<����h��Ο��	�L�IN�R��B�a�0��A����-�I�����	�p�	ßH�	ӟ��%��h	�+[*������ơ:8|�IٟP�	ן�	������D�I�$�ɚ'���R�P�EB�D�w��*���	��p����I��t��՟�I� ��5<� ��QgҞ�ꥂF�՝a�����ԟ�������ϟ\�I�X�޴�?��H����%#{�$h+𨅮ZH
��Z�H��cy���OڝyC��<�&prQ�I;�D�xJ�|V�=�3����ٴ�?�v��j��<���5���p�X lcd \���h�7��l��h�Z������	60�Ăg������-�M�o�H�B�蛢"�� �	�<�6�C�T#�x"*O��' Fr���ܪ�gċ��yb2eV�)8p�M�8j����<��'[|�|�'�6=�f|zv.	]���wF�&k�t�wa�O����F��`�	81>aKԝ?9��
��S2�΢F�l�#�a]��H!�A!J��' ����TП�pa`� ��de�@#��-�JX�	<\m�l1�+�(�ޱ�r�A4,��VyҞ|bAQ���ٲ�yR�X�i�l��5K�vj��3Â�6e$������n}��'��˹c�t���/C:�C\?_�\������q�KC4�y�Np�:��$E2"����GP>	�*�O�L`���>Z�� 7iH7�$��!FzVԌ�-O���W������9O�˓q�0�Is�Y%6��H(�����+d�3PCa~��{�J�D�#�1��5HEoF&]ؒ!�Tg�%'�T}��.��<�Z���)�O�]�"�ٍ��]�J�<u�mh�����k�
�y�n����=d��eƓ�'@�u e��<��'r���Q67#�	]�4��|��}���k��9֪�!
IH�'i� �Yeg�b���S7�d�_#Jy�&d��0�F�j=l����O8�$Xn�n���U|�����?��o=��	'A�1�~H�v΋A�.�pϒ�6��6m�O�ޅR3��O�ZѮJV}��P����?�l�T��+&���p��\ H*����vy"S��%��dK S���5#��8�$#�"�N#UGL"k�扡�MS�W��,���'���'Ì��B X�9�|�c��V+B��n�q�A��t��qI�� ��Ȃ�4���]�T/z���?O|�]�k�T:9}���."Ŕ0��5}�r�K�	P$�U,O�ԟ.Y���'~�)aG�ς{�N�� �˦�c����pb�x�!����4�?)�K��<e�G$v⠄B��ʀM����[�ʡa�'�ơdA��?ͧ2K��Xw^b\=O\�l� 8��љsڄ�i ۿ8F��'Jn�ɐ,�<�'�ݐu��Ei�������Th��e�4�[�����po�p%����N?%c����,�P�2�N��b-Q"D��/f�`"�m.?�T�`������!��0�?���ğ|E��I�dTtMЅɗ�LuÇ�L��H�ڴ4��A� ݺm����uWč;�?I��Z1�.)D,!�̤Y�i�2�ɨz�� �}^�!DV�<!��|Z���?1+O<�(fO�0$���{P-C�@"b@��9AT��Sk�O0�$����1Y�����ɩ�MS��Hw�%kai��%�z��sfב9'�F��+B	�G��r���᪐ʟhG͐H��ܣ._x)��'`�e�e@��u@֜�7�3	��uϓ!j��}�ڬ���'Q��'q��-�p��0َ����xI�]�Rkk*�)a�J�doRa�	��`�I�?- ��Gy�Mz����<!K'�Ys���d̨^���nڋ�MKCOA?����'cH��]w��	3pbʦ%T��bի(7NTBt �w��"0����_-�YER����oٔ����.�?)��!V��İ��N C�~qh���?���?�����d�&j��xa�.�O>���O@ ��K%�}�u��7��O�#����O��mZ��M냥�j?1�	_*}�
��Q�.R�ѩO>vT�[� �ٟ4�����|R��`7f��X,����`�ןP��jТN��P(�#j7�����ŋf[Ή21�'���'�dx��K ��O���'�2��F�=�WO	?E�r��7��[�d��7��ÄY�l[۴�?�O�W~�wN�)
�*'}�`]S��Ңpxc�D�>M҈��
w�(]JUNK&E�*�����b���{҈y�U�ŉ��z��Q��&�`׆�y�I�th^vy���OT� Â�D���D�O����J�   ��<p�@�\)~t��@��O,=��ʓU�H��ԡ�?)��?1��U,6��'�?q�b�)6h !§��0�� �23(�	��M[s�i ���'Nbݻ��(�B�'�+
�XE�k��B<I`3���̐�\�<q`�ܻ)��$J#!\���'���L�'�̕���<f\��`�~�@ $+�6���O����O����<A�C1h<d*��J�E�԰�$�0 �P��`�R,�6�'�pxc�OX��'�x6-\�EH2�	
w��b�W�\�Rg\5Q�Vx���	W6��n�u]�I�L�u��N�?�9H/����=� (�JF�ڶ9kwnޛ01���AT�f�l�O����OF�i��.�ؓ��N҄n�D-P/-����+Ř?�"˓�?	t��܅�'�?Iзi���I��y�#�6
4<,#1��9F!z��ǹl2���'���a&?��O�.=ҿ�^0��-n�� 3�B#}�If��UD��РEl��'���{4��<�7�'��]9��]�I�2�'��b>�zx�@�9A����#�'0�I ����G�،��͟X���?�����vِ�����/(��K!�->l�T�I̟�o�:-�h�	=XR(Z�=������ȓ-3�@j��k D\����#I���%�$: �t2O�t��?i#-�i�	�S��yP�Q���&eoRY��*����j2�?I��|��?�/O��� �8oZ4�2 � nÄx��,0$Y>9Ӵ(�<1��it2(4��ĉGy��io:�qe��*�Q��#��`���s�"����_���C�M�c���$E�/hKZww�ę���<1�WY(�@���(F�F5m�PH��$�?A���,b�^����?i����'&ϓ����%<��J2gY�Q	�AFC&����ID6CH@���O|���P`Qg�<�մ�y`O�Ah�LI�ٸGA����M)8��6Q٦U[V츟�3��J]���"������%*w+Κ$��}� �S�?VLܚ��@�y�,�pD6���+\_�ܹ)O>0�	�}��y��������O��]�:0����D�Xy��@�������	Zy"��=� ���'i��'$��i�+R�x��T#4�T<����'��J�Oh��'�7�Ц��ၷ��C0�߬b
�IBFB6(�¥ܢl��j�<O*��@ݗ"z,6���<~[��$_�-"I���R��@<`4�	��?����?�/��B�d�K~R��?)��(�BXcs�R+Tp����̖�,c>-����Ti3�d�/��$�����I���Ӽc��^�x&���I���� Vzt����7)��DٳCQ�eX��iA��ݟ( w�P�U�.; �:�Qb�%0���Rm[�Mx��W������pBcK:/sJ��Iǟ����?y�PoS!YgH0���]�2���g��7�(�'�<���@�I���'��Ov�-��]��z�%IJr ���@��~�qb�^�����Φ%9ٴ6M<L�.�)p�$��?��S��L�����B[Ƒ�pIY�z�<T����-T}�e%q��q�	�<��A�7zqn˓K����� H8,�=z���kA�(
�<�6�V�yB�')��'��_���cE�,���4,h4-R�L�i{��I�]�֐���M�) t��'���?�شm[�3(�"1�H�����~G$,�/2��;� ��w����:"��s�v�- p�J�p��$c�}S��96���X��%�v�G*E��ݣ*;%C���?����b�Cް����*ۭ+����-�6"^Mk���6�?���?��@p����'�?���ip��S��y"*�
.��"4lS7��T��t���'���Kr�|U[��|�� J��u7#�=/󤔓]�8
$$��s���cC_��ϋ��?��FQH��I �?1&�E�E褰��?a����y���ݺ�*x9�ߓf�$|���?�)O="X/o����O��d��X�@�lW�~�nP��+��FU�]YaXb��I��dTЦmkٴ��}��#ؔቆ�v>���
d`�V�؄%W��0���2)��jͧk��Ѹ�/`����L�R-S�4�Z�L��$�LùN�V��� Vz�l,J��'S������'��Ok��'6�I?+�P*�� ��
[�ȋ*L�$l"7h�>A��'.87-�O��՞���,OV6ڇ�(8�(ٕM�H����l�ml���49G�3K�t���x�l	a�͵)����	�D��'p.�`��-0����8H�������(��x	nD;@�'H"�'�T�Լf���	"(Q���]�f�9�����O�%\@�	ş0�	�?��gǅay��n��n�#v'ܑk!*r�AL:�L���l�99ߴL�<���	�@2��k��u��;_Ζ���� s���3ӈv�P���<O�7`�>�?�/��	��?�⎐t�R����ԼP� IB���M�WH�1ɤ�����?y���?�*O���#M�
8��$�O>�$Q65"f�� ��i��(ܫ~�����F�I����CӦ���4C�F���v@�Q!�*(�`'�M9a�:Yr�������#:�,��C7R(E�k�|���̟,I͊=	Ul�ɱlՙ�"0�7gT�@� #�'���'W����	l�On��'V�/�85�B�CA`]�Nbh��ś�����L`f���T��i�4�?1֫�y~�w"���-�<pJXK���2_j�Xc �I����d� �c��i��]�e͓C���cG{�E�Q���2��=�T㟽Jw���b���1��4Cf_� ��y
t��/��?1��?���6.���֝1��H�����HZ�CB�Ĥ��D�0J2�H�i�O����O���C�D25⑉��_�����蕨I��82T��Q�4	���IT�~R׶`�P��'�ҲA��m���f�M� �$*Q�B*<h���>g/�(�M{"ݙ�B�O�`{$H�xy�h�OP�ڠ�W�	@Iz�J�r�j�IG;��t>O����O����O8� C� ;���6�?�%� =������;:B :�ڹ�?�i��˕�����}¥uӎ5oگ 8F�B�͡xp�ǂ>QX�:T�0Rڨ��
P�K:ʴ�	�0m\�;����ra]�yr����-��+\��d��N�c�>��U���R M�	蟤���?��g@T�s�!��]�F��p��+	��0����8�	ԟx�.2K^�ӟP��4�?�Ī�<9��,5�R����.�p��c���g����Bd��RBb���M��'�4xj\wO���c	�O��93˞�d���ȖHJ�n2v`�e(����+�`"&pk�W��A�kP�0��-�?A���?�a@nr	ׄl�3���%��y���?i(O�J$j�L ��O����)�e�2}���k�@�N�-��]�h\�I���$�O�7-�?O��H  ʩ�O�n�s��?$��1J'Qu
�X!BL�Gn5�A�_�M�$�Q����aV�0���E�����9{e�k��H�~����7"��~�\l�	�<Κ�cŎΟL�i>��I��'��͒5 ������EFH�N2��)��e��Y�_��r�4�?�F�]u~�C�>�w�i������,7a�7u��M{�z�21;e&4���v��+����U�_g�9^wŎ=���<� ~p�đw
�b��-h���{"�'����(/�"4�'��O�d�Ox���S��˧x��5���ֺX�rArt���4"��5���������?)���2ĢQ���$̦�'"�V�z�霐}�Vm;P��:{���;�4i����!�~BI o.��Oen|ڣ��&��q-,�&�;�b"�Fu��"
���9N6z]R��'66	�W�<b�'p��E̝%�R*W=4J��ȦI6Js����2�'���'��ɏ{�\���NNß �I�����E� r��|�fĹ*�XZdg�럌QB�%?��X��I���3Pe��?q�3k��|*��8u.�3�����C`����x�юBa�$NP�;:@<�O�(;�&p�m8� �"pMNe1a�B��iz��ƓQ������?i���(��$-��䧆?��?qa�4+I���8_i|��q����?�`�9ɂ����?1%�iE���4�d�B�#r�h LT2d�8gJ��3�,�����䦝s��WEKB�;)ةhKқ`�4����@<S8n�#o�
.L�HW�Ð]��%�\�5��+'P�����l���ĭ�?����?i��XC�������y��bڡua��2 &���$O v<�� 7��O���On�ɍ�`Pʓa�:���j�����7��T��bӒ��D�Ҧy�۴Hq�|����.3z���1_�eA5���|mk'ˎ�Z'�2�j��Ѷr� }�tc �uG��6�	&.����;A��e�/U�TE��7��0��@	���J���'�R�'��[�����vڵ�I�*����!��F�
yr#7/`��I��M���-����'�~�m���k�JU�礏�;?6e#�/�8�f0��ʚ�ow�5"��M���:X��-ԅD��uW�
�O��y��!���_�F�yGcS�v���I���$"��ٱ��w�J�A��?	��Z5�I-�����K���y���cϼ���Y0�?����?94.��T�v��.O�m���K��i��Ȧ��9V�<���I� ��yl�:�I�<j"�b��⦭��$-��;	�1jD�'4���A9V��P��*B�yd*����¹b62��I�%�<	�'�,��1�'��a�N:l "�'wr�Ǡ
<X+��:����׭�Bh��'��I��XM�"��ޟ��I�\�Sw8Ph�B(ܙtA�PVJ�da�ź�A1?I�\�ĉ�4MY�6&��~��P-zH"��#���P��^Ug�1��^�.D�-۠Vz`]�r&܎W���͓��}�6��O�Epgo��<���n�
�	ҤNy��%[�膫��P���g~|�g���?	��|
��?i(O"YS��E�jܠ�q#Ö�9߰y�o�!7M��*�H�<ᢱi�r������Gy��i�u+�/��@�6�b�J��D�T�R�p�P�)��I;O�H@w��0@0���_	i�.aX]w�Kd(��<�r)\�7Ѩ��Qp�t��q�:����)�>u��	�?����?��'Q�:d�+����BB5&�d��L/G�q���s��C�O����O����_�ʓ��w��܋��A�+W�E
c � o�q�1J�O6m
�c��D��B�ơ�7�O��H�:t뎌�(F +��׉X�|���Cˉ^�Zl��l{���%Y5rΎ&���I�.�~L���4m�����hAǤԧ^�L��-Jw���h+�şp�	�h�	\y)�(�у�'w��'�H��'n�H1L uO�u��)��'i�u��Oʠ�')�7-NȦ�SF������ҥ-^�DHs�K�4�>	P�H�)O�`�74O���`�@�h�0�:�O�k���4x@���O�V=�v���/~��P�۽/z���g	���O8��E�n&^�P�!*�	�O��d�O����zƺq��. <�|C$`�OFMP�g_�J2�ʓCg�&�'b,Q��O�.��6�~Y�f���E���%�+(�ҩu/�6��l�?`�$8�C�ĺ�Ń�%�y�Ϝ�*aŵ��ѐBřP�b �~�p���I(h���' p�'��k�f�56��'B"�O,T����7�*��7��#�
��Ć$��ɿh�n��'�۟��	����S�
Z���'b �s��Z�Ѝ���E:3Qaz�.�>��i�T6�J�+�����$�SK?�s��L\�}Õ�çP�9a�Y9M�yD�RaZ�Z�M�ԙC��L�)�g8O�����O� �F�2p�.�c$E4p���25�|�0���O�$�O\�D�O˓DI�S��?��!E�'l� �E_�=�N�PŤ��<5�i�b!Q����Iyb�'C����r�ND
�ΞY��*��L�H�6&��u:T
@'&1�x��m�B
t��3�&%2#�O�h���w/u��d##�P�:����y�x�E� BN�͚S�'o��'
�$E�R���y��� A�b�2@��/o� ����t���'��w��(�X�p����oZ�K�j���Q�o-s��#ώaE�\��坏�~���*a��ʵ�i��K���Nň/���I�f�V�pvf߬Ay� �샋 K� � ًga�'�2I.��ɊPl��I���)���̟8��͟�K`QT��c���J#DQr�E� �Iyy�M���z%�'�R�'������`k�����:Y� $�9^d@��O�d�'�b6� Ѧ�S �`&%��u���ۃ)� ɳA�3F��kE�,c ��q�͸5�21Kt́ N�D��)�k�F���qt>O�
����E�yB؄��%Q+Da����?f�b�j ��OZ�4�����O��R8Fa��9]<��{E�ħ"����Ӷ�q;�BnyBLu����1G%�	��xӀA��
�L��LI@N���vehVi�Ŧ���@!Q�i!��HZ�<�	,Havm������P��y��#U�:�H�A����4�Ʒv�1�R�'����q�/i�R�'���O��� Y>	�)B�a�T�B�e:,���B��~o@9��E��<�	ʟ(���B�j��'�r6=��0��+�B(F-+$,��r،��d�¦�b�4R���l�ċ7(��?��S/W�Xs�i��m��cYS y��E�~��3!�f�̹b��:\r^�t�V�+v�I(%$��*��Hџ�{��-M2dxҀ�> � @:������Ο���myR�Vy�Be�'���'�(�r�����𡓔H�u��`��'����O6��'��6�F���l���A ��3?���!L�օA�g�Y@B�x��O�-���\~"��@�6l��d�!Lx���Y0ڔi�~Rl*�-����:�:g����O��$��nxd�k��9���O^�$�O��J1��@*����'Ma��r�i�O�y@A��a��%����'����O��u�t`5ǝ�a�P�f�]5�j���y��tmڋ_�dA��?����{����K<*l���;ƀ �q�1D�=UB���b��Q\�<��R�7�A��n���/p�*�KԠ�OP��O��I�����
Mo`��3��P4jĮ<ᓅ	�I�	����?	����I1����8r�@��o�� !��H4 P�'R:6��Ц	!G����#I
���i៞� ��F��4�@69��%:�*_1#�D�A��Ff��ތR���F[����8O��X���O�ڕL=	�t���, 8:�|�V��P��}����Or���O,�D�OD�3�X�S�?�QER"%�p=���C�$i8�8����<Yf�i��A����d�|y��'�V�J$FU�A��E }˨�;r"�'��t��-�]Y�4�"�X�7"IFIK�Y��,��Zѧ`��rҁ���s����
+�I1�88Ș,��$S�����ݟ8���d�ӳYy�%?睌����3\;Od�-���5S���Iʟ��I#]�f�qc(�LyRFs��$���ּ-����#]H�������d���O��R#,Q0vq�6-���4�h%T�ȟ��?���/bИа��K&#����G��&�e�C�i@R�ŁzI2�p���l�P4�'��'��dh1ɕ�1�D���o�R��y���'�I-� -�q�q�4�	̟ ��)SH��5Lk�E��@�Yg��;��>� Y����M�E��?��	��*���ӦPi�hH�D=n�&�B$�Ŋ5.�IzB��4q!.�����m���6I2��'ݜ҂���ytcP�!kH`ytF��Z���DŎ.�?!g
�I�tݠ��?�'�?y���d�(V�0cFa|���"��8Ⲭ�G!J'��	�M��|�<9�'�$�l����5S#>9�B/��-�h�!�3^�"7-M'�"mK#�D�~!��q�OBd�M�u�Ǜ�kX
����0CaD�gUЁ�4�d3u���.��):�x5��'-"�'�����.���5WfI�'�dkp�PK�l*m����E�
��蟔�	�?U�6O.?!ս�y7HV$<У��D*�Fp��ăI�l7͏Ʀ�*Q6�?!@KĜ9.��'*9��!��ȳ`���B��=u��I�?;�ó��<�Q�Έ-����<\�4�'ܺ� W��$��O��[��: BR�|f�s�M�"�'��'}�;m���rj1?!��"۾��S�ɳz��]SJG&:�X���'D�\�VM|�B�� ��ȟ���C�4S�ȁQ�G�`YԘ�����z*a�� �O̬��b��A���Z@Q�̓�ug���?�wЌn�؁�
�9��(�ׄع� \��a�Ob�$�O:��V�I5Gd�����O����T4��#��X`�
᠗M�)Iz�d׷�8����<ᡵi���͗��4� ̉b�bGDM�w�4���	@F�l�GDĦݒf�8w$@,�e�fH:�	�T���s���PYS�L�m@�B%$c�T9���Nt�+Or���,D�2<ɶ�@ǟ���������2�bɡ#�[�|�ЭE4m34�r��Sy2F+I�e�e�'M2�'����j���8I�t��+X2���c�+�Ҭ��O�m��M{�!p?����'p��H���?-���V� h�:�+��iM�*ب{�T� �D�D�2��W���i���O@��"Dy�)�O�h�#�R� S��7Y��
"�$j$HD�B/�Of��O��$�OB�.�����I��?�2.�VU�	٧A��t9�Q���<i�i�R�����TU}R(v���l�p�@�y��ѮW��ҳc�P<�ݐ��N�^��*�*D�@S��	�"���q�����"�C��)Q���j��P�� EA� i�1�W�˅J����\-f��'���O6r�d���w���`�O��zf>y OHKNP�'�'���'���c@�>�剻�M��Vk���I��͋!��(Q"&� G�h��.N?C�&K\3��|
%dV1V#&l�GLC�<���<R>"�IwLr{�Q���W_�!����O��y�oyrG�O�H��U�Eh���O^��;k�y��"^�o@��fNݩvZ��$�O��S��x�d������O��i%X�@����K�>�Q�M�&#���+���\ʫO؝o��M�"��T?���Q&/��S�UB��@���RɄٺ��]KW�`"�"N&4*U#Ō�:�����{(˟$�4�����*Yƨ��#nކ؈�[v�jP�	�h|�$�t��џ��i>��ݟ,�'�<�y�͓�Y�d�Z�@�4��px��۸Apt�O4Dm�ϟ�H�(9?�TU�4SشL�N�A�\�)�ǚ�\G���iR��G�U��:|)b�ٲPy��Z�~Q��;|�!�"~���/�6�L!��#�բk�O<��-K<37/������՟|���Pn��O�qa���_�t�Cb	ԾXW�E�P�.�*�'���'���H"����զ��=<��y�� +�z�y�T!9zQ�۴]̛���-?u�$��b�p���O���Gý\�� �O٬QI�zR�9PѬ-��ɣCK����'�Nm�2I�����G8��$�� �󧍒9$��ɝ#�H����~`�Ȅ�Į)��������	ǟ��'��Ir�	�/�'%oOC�|@�������`�[�b(����^}bdmӸ�m�-l���I� ,*��2D���X[�U�}/�,����|��DϧC�
��"��"����w^>����O���0��'/#�I���C�����A�i@ �����?9�C3��'E��'�?���?��E'=OP�:���&[�����P��?�1��
'��@�-O`xm�͟�Auh1?ͻBe�]b���&q�9�΁�9���+$��@�Z0�iq�+�gɆ|�ȈS���.:2�A�Bj�9����ϲt�\iSdmJNĪ��
�(gg,�+O��Ɇ;�r�Y�&��������4��<`��
ɆTQ��Z�� 4 R��d�`yr�D�E���'�r�'����͕���4y�az��K�P;̅A�V�2���'�6�ئ�ba䳟�x�/O�(�~�I��p�kU'΅z����l؃K�`x	u��O��X�W�ԍi��Ʊ9X�ۜ'Fڭ�EV��b��&��T��	Gh�-�c��%%_($.�b&�@��h��ڟ��Iןܗ''���&�NY���2L��R�B.B���DX2Kt����Ú9�������ڦ�"ٴ-�Љ+C�N{ܖ��w@\�oq� ��͸%)�p�WM ��ܪ4� �jq�NI�b`��ȟ'��.���3�ٺNN899�ߙXIF��S���xj�S�k�۟�	����"�-�9�Fq*UgQ:����<AT�����OJ��O|q;5 �}j���O��o��S
{�4چ'�
5,�0�D۬a<�m�Η#m��	>P�x��cЦ�S�uRh�8����"�	�&��� �$J�g%�.\��+s�&�����y�����	0�?��oL�/��4����?���D��,�CdY1R������)~Z�L����?�,O`٩��2����?���Z��z��C�>��s,L'�Z��Fmk~2o�>�P�i�7��L����6vZ����O�6H�`�"��e�剢:7����
xN�!o�8m��R�'��n�g��	g��
��$��)�?B\�a; �O+D��Lb�'dZ�����:�������'\RZ���c��SN��c��$�\�C���z Ľi��PQyb�n�z�d�p�����d��ݙ��W���d.\�0Ed(�b���M��.���K��� ]��t����	|�!����M�G�i�`�߬A����e��z��a�O�Lb1�H"Wv����O:�d��������|�ӁF:<�vԫt4��<��,��1�ٰVaϙ�?Q��?��'�d��,O�!oz��`��&x�����G>`�U��h���M�Ѵi��1A�'W$H�O������W?��b4����&��W�H �Ɯ�iv�Ba���<�]j���׎1��'�8�$�#R�Ę���O��Q��3X�@%�����Q61� .�O0��O"�$�<�2�y$dp�,O��d��e�����yXh�`c��w,Z��	zR��K��	!�M��i�2� �'�<��W聱w|�Xpa[)l� �@-D�����nA��kÁ�B�¥d��<�Yw����%�RD'�!�^�×ϙ�LYq��Թ)͂���O����2�<��b%���OL�4���7c�>^icS@�g *��O�]ÀMG�v��I��M��=7��y'�4A�8�aI�,+_�1a�a��<22	3�G84M�6́<k�t@�&E/h߰i��O�|[����u�k�b0���a�QT���O���!V�\wyҤ�O��ԩؾ'\���O$�����q85��3H�`�9�ώC�PQ�v��80Y�������<9���?����d�'���n�JTp�q�  ~l�X���>�ûi6�L�P�@0�ɓKg��R�?�"�W'[�<��N��X)�L�ݺ�����!_��6V-&����'v�pȼ<a��'j!Ara^���-X�Gό5�!��/ �U |�u�'+"�'�r�'��b`J` &f�4��#H)TM\� �/^=#w�6�f��`ݴ�?!V.�i~�
�>!c�i�7�.��е�T�b�(6���H���C1��&~��%��oޛT�Z���jR���]w�|"1H�<�]w����HD��e��I��	�;1ѕ�̇1Z�����?9���B	X
����CAI���6iYi�r�k�-�<���?�dkN#'�$��'Y.7��O�P�5Ot�IbZ����j�naY�K��gϤe�ɂP��jV��֦5�S�� ̂!j��_����	 }6+4O_�w����B�5gv
A�@.�@�"�)[��c�r��>����'D�'�|dABK�&F������@t`j`�'��_��@L�u�I������?IJs%]/D�F�ܣFuX�s���*�����Iԟ0n�PN�@�3^q�m�?����ޚ(�x����H?{���[ĉ�_���M~�����`��;lLD�I/��T�.O�}!c
�!B<�9�L+(��,c��SӟpA$	Ǟ`^�	����ٟ��	ny2I0Ft�Hse �;�ʙ �&�!`�LqU��Ibb�'�Z7��O���v���I�OF�m�r���Q�B�0�!��AҦY���uӊ,C���f�P�����v�h�D��1�Yw1p��H��<����~�p�;cf�,=0Pp��韄��w�n��rC�0�?9���?��'?��p�)�D�Q�?}�~���K�:�&�C��&�n勠m�O��D�OT����:M~˓M盞w�¹��(�]�x�1v�P�G�,�|�\�oZ�^���	�{r�	IE�����Ĩz�z8Y掁39��$2
U�v���ڙ$���)D<Oڨ��"��y�	=��I5�?�W�i�AiR��Of��U��	�J��C*�A|�CP�O���O��$�<!�	��*�X)���?	��
Q~@���)@�$����̲u���s����'�����v����OB�҂��������!�h���R�a��R�fM�@�'!�.QZ�p�!�C�Z����u�b��y���Rށ����LcT)��LT*e?�Y� +�O@���O �I�Ǟ)؀��^��O�N�! zb8���l#L,�ef��l���d�85�jٻS��<#�i}b+�/��4� ����(*enD��*�	D5(����%wŘ����Ħ�(�$�G�΍��ŝ�]�I% �)�����·����ǘ�B�K>Cn���������3�� (P�`�IП��I�?����\�̥;P!R�E�Xj�'ѿYW�ؖ'��]V^���?���r��h~�ʄ�W}l�F&`��5:d��%D�E3���}�:=c��ȟ$K�LE�av"�I��ڌ!0�F<,�D�JP�	k 	�8,�$Љ�(X6���*xl����a��єS�L��y�����8EOT���C�5z�zr�@�b�XP���?���?����&�x�9O�(��#�h��q1�I�FsB� 1OPhm��|;��9?�U��!ݴ@8�F+N��xa�b����j���`yǀ-����A���MA)7U�ͬ�f�N�8 �T�;H���rD�DCc!uB+��h9�+�
����G�ΟD����T��8�pl%?�]&x�R��tᅸi�5�Gą�~
��?1f�A)��%�'jb6-�Oh�!9O���1D*jЂ�`�#p�Yf��E@��Ɏ7�蜱v�Ц���	3�(2n��'��!�\�o��(v��'�"@�V��*Rµ�I�y'U�,OVQ�	 Q���p/P���I�p櫄?2T,�SJ�E���@D�WߟL�ISyR��5�"䈙'K��'0�T�Ĳ"�¼:f$Pu��`�*).�ڠc�Op��'��6-P٦5t��?�vK�˚��Ybd9BW*�*}n�H�(�+�j���i֎b�4��D�',P��韚�	��'n�}��J�<��l��x����:�z�IM�#�¥ّS��1�'��O��'��I�X�m�cG�u���@�#,<9`ĦA$�����'Ϛ|��O
a�'O�6�&]HТ��	}�H�J��ݦa:��Qi�*�I�ݵ���I$!�`���)���y��i�*���ǎ J�F��?i1�'�&4��\@:"�'�b�OF�ș�U>}��KےO��˴LAa�d�w�ل�f��e�e� ��ӟx�Sj��g�wʹ0�t��7:�5�$� �(p��"kӮ�mZ�A �#��_a|���>B8�kjZK�? �ɛ� _�h��nټ���a2O�9bg	�?1P$ʹ
V剣�?����:(,ft���;��u[C�߯CI��ã��{5@9{��?����?I.O����G�~����O��D0X��84G��pش1"�h�|ˮ��"g��������Pٴh��A���'��!VϳJ	V|11	En�Ժ�dۦ>}
�Γ���X�&E�.J���W�	[��mY��?�f�7=3��G(�<nXE��
k����OP���O�@�%�!�����$�O���Ҧq`�5CPf��f�ؐ���_3<�DS�'aK������q�	�w!��Ӽ{08^��\��A[�5��s��ͅD~�&
k���F�g<9�BB��_x s6�'-��q�d�غQ��>Yx,�y紨���.R� hpN_br���?qf�˖}6j\���?!���%��hi;d>����
�(;���+O�|R�kQ=D|�ʓ�?��'��,��J��oW0��bf�����A���	��M+��i;�а�'��r�<�z�'s������8BZ���̀�:����B+��?>!X���<���&:�:���/u�Pt�'d��$U=9�$1��P���&R�e3�DЩZG	h���O��d�O$�D�<��̒@ ���XvX
a%@�j�����ỈP��͓RR���'$U��OZX�'2,7-�т����41)SVf]�n\2�Y�ʪ9A�d+��9���Z�p��!Yz��Yw��`{`ΐ�<1_w�6��Ю1X4B�E�8p�Y*f%��B�X�#`�E3k�����O.����ּ�p:�9�>I�V��$1��ńA$
�P8j���O���O�����`�>�f��'�d�8�'� y��.� ���{�%��
�hH�HP��~�mX�N�ry�u�i��T�������`Q���HK
?Ьv
W;gX�1#5�ɧJ.T;c����[��ã��͟����j�"���՟����Z��JVD#.�b�'�ѻo� ���T�'��!�Sڤ6��������U��ihQ:-m&]���j��(�=?�bP���Iʦ�â���<�ԯ)+����36KH5��c_�{�������|L۠��d�as���2��g��B���O�c��by��V1yO�$��+ˎΥ����$����S.k�8��qK�O��4���$�OH�|�$(aT'��^ΥA�Hɪ51��k�M/dӊ)K)O��l�џ�"��'?9S��l��9��� �J�<^���&�9Z�f�۴FlQ�v�%C��T-�<iY��� ����͇"�y�K�v�p�8�E���p�Ś�?�0�'JAГ���O��'���O��IA�V>�`�Ç�Q
��``!.+�$��$�p8U"FHMΟ��	����S#Ԟ��'<6=�f=H�'Ҿ\|=��ϖ�R"r�g�æ��ߴ^Έ��5 ���%%�e�E
�܄���37|T�4NQJ�f4�cC)q͓H^�r��f�ȘB�Cgyҧ�O�a eG�$H���D��!�ڑj�@�# � �p!G�LV���O����O��Z���y�����?���?U,Z-D*� �a(��pv�E ��V��?sMK~���>a�it7Mܝj���YMV��(��))7�	*�|�б���y"�N�0�6�I�G�\�p)�-�<1҄6O�d�4lH�<)������]\hqyU�V�Ql����(��%V[���d X���D��՟�`��B�T��LF���X|f�$�	��ă��O��D�)�I���Ӽ���%1��i('&|�<87P$X��<AG@P�bs��/Z� ���6(	�e�z�'��
�Oắ1-j�3�:f����" �=�C&W���ϟ�
�DYt~`���ӟ��I�?ũ� h��}kv�5ny�VgΦ+ٕ'$��I�B!)�B�'��O��Ou"m���D�cSJ�	2q��kċ��Z>��?Q޴_u�]��=vԹ3���?-��<��,Y�*31��; "K?YW]�p��U��|��Ee��kQh2��}��B��+���!�J �D��
�#I�:����-9���'q�'r^��( �<_ĸ�Ʉv���aF�	^�@$Q��S:��I?�M��&�E�'u��|%��"`�0�k�\4k�����V:>T(Ya�_~Vy34���Uoh��Т�O����5�u7
1H1��ϓ�uh��$#ܶR�B(���<�(@p"��Rz�!5����?Q��?�'C��D�K~λ��	K�Ä�yజ�D*�PIf����?���m��x������d��q�	)*i:�	%f=�a��N���XQ�	�/V^]j&๟x�Ώ�;ߨxmz>��%��"�T��t�}�D���Άl0P���
4AA��!P  �6O$�����<�'�'|���'M��'bȎGj�8PT��5eL9��D͙�r�'��	 #M����~�p�	۟<�SH��0p�
Z�Y���g�h�6	�q�??�'U���4f��(�p���IP�L�a�O�:����_	$���0��V^r=�"���[��Y���_n� 8��Jb��柘 r/N���V/Xx>�p0�1l���r�s]n��Ɇc,�ң����i>��	ߟ̖'�8)��Z�Z"��7n�$�R�3���� 4�RR�i�4�?i�k\@~�,�>i��iC�U���R��U��n��S (5q4�{�P�u+�� ��)
�"�$66��`����^w�p,�E��<9� ۂ��iEN�����g~����d@`��ZLd�	�|���?������x�+T
�p�H��J�#�n A��28���������?Yx� �Pyb�d��ߥvº�86��:L������- �PnZ�M�9�"�5a�G�?�Ӱ:b�q���8��3��.㦀���P4=8BuRů~��"C��!I5�k�-剔�?9V�F�n��q�mEc����<�ZD
!NU�$�xq����?���?!+O�	���x�x�d�O��D�,� ���B�x���䇅�2����)�	)���XǦY��4wƂM��j�Lp�̌�=Ϩ�K�[�fdLC���h�J��:K��p��L�T�(&Ƚ|:Q�ğ䛲���Ľi%�ݧHN�Xi���k�XL*f�'(��'*x<���0��Op��'��'�7�9�-B6r����[�]vr�#��1��'�r�j�B��	/EF�i�u���Bs2����A�&Ò8�,W���1�D�˾�MƄ�%���3��ɒ.�͓c����`*y��
�B!c�k�#^�J� �=02��B�BJy"�O��%�
	~���O��d�:(´Ɨ-?�x��fƭl�^0���%��˓?��d ��&�?i���?���2Y��!*O��ya��:@��&ԭ߅ǽ9����'�7-��)��i����$���� �� �m��[�����FY>!Ll��h�&,Tݢ�9O�a�򍇶�?�(\�H��	�?!��޸[v `��	w��%�$B_�I���#���?���?���?Q(O(9(@f�>kF�d�!O��`�Y8�Z���c[�$����	�O4z�x��	矜mB[Җ.>o�����	�� &Hա9Wʩa��>p
=����O���`e�=�u���`kFa̓�u�*�ﺸ ��ŉ[�|�G�/{y\�S.G%W�^�DE�Od���O����+ ����N#H��:��J9MB0D�Q�؉Dd�d�O���J?@;bq(WI�<��iT����yRK��d����I^MA`�*_�Ј3�'3����U�e4��O$�V�?�x80d�'�r��CHݠEz3
f%F/L0[u�����'��sb*�<��'�Ҍ��Y��R�'5��7��XQa� �^m�)�E��:R"�'d�	�m)�I�D�t���	ٟ4���0��h�eo̝H�T�9T`��N��(1 1?�7X��
�4-���gґI�����C¬���OY�Q{wb��'yh�ʳ�K1nbA��fJ
w_��a��&s���ژ'f�.O��� 
e�ʓw��ɱd�+.�аⰨY7^��ib�'J&�4ѯ
�������'��Y����Ʊ|Ad�a�/�Y��U�e�@Is�����'?�v�i]�������l},dӌ�.]���� `=� 
o����6��RzYj�Ϧ.��A9���O�}�� ���u��ϓrלyΓ�rQ��d �BD��	T&6�����
ڴ|_�ź��[��?���?a�'A�`H�+�*Z�b�Td��%�(�h�&[
(�p�ȁ<O<���O$���\��	��MϻM|�Thv(�?:\�1))',.��im7��pH�ɿ0�\��K��~��N�M�����(��D�VmR�c���D>O� �ҡ��?�a(�V�剸�?��(D=x4����9��av�_20Ų����v�@���?����?�*Of- ����B�����OB��W�$S��V�΄�F�F�.����'a`E��O��'d7�X٦]�!����[�I$h�,=)�l�E^D1 S'n���ɱ5O�%3��PiT�q��E���S�M����62u,Q��C�3
���RV+�*t�hP*��?I��y���}N�{K~����?�;p	2�@6𹒵kC!�*xK��A&P,���U ���ަ)���>$f�Ӽ�!��**�\X�����dd��Bj�	9XiC�Ε2Ji�V�½�
A��g�	{��H �'�|����庯1/v�ܡ"&����L'04�E��Cۭ��Ā쟔����'����ʟ��I�?�`�k�cDX�GM�� �_f+NF���$�'B?������O`��O��)�?o��)�O��3@��L� �x��b����Zy})e�	oZ?�d�	z�x��th�Z��B��x]�2	�|lt��V蟑;L����.�z��6O�(5+��y�U��	�?�BC�Xt.����J'A�<�,�]�	h�
�?���?)���?1+O@����Vj�d�T�V�`D.4rJ�X�H�9K��D����5<g��Q��Iޟ�o�b~�UR����S?����n�9o���3$�� D��8�,ԽU�N��9N�1Z�� 33����Ɏ�߅�R�� �+�/�5E�j�qG��	��c����	��|�Sf�%'?�]4W�\MрF�5[.�8�  �2-@U�I՟x�ɀ769�/j>Q���M��Z� h��@����ϭ :���u��>"�juɡ�X\?��Q�>����|��R�#;��`��<��AދxX4���ťEbZ"��7X'��Z��c�\cVDy��O���!b�0[|���O��$�*�P/Q}�ac"�Rì(a�'QbT�<҃*�U�	П��I�?ݡ��/-����C�8b\[7�Ө�.�s���M�i{:0`�'Nź�i��|��E+��� 6d
8�ipB�)C��r����A�%!���韤Hۄ>O*|{'*�<ie&L�/zU�բ�\�P*���.�lAEe
H��'��O���'�削&	��s���{Ѻ!(��Q3j�DI�2
�lA�'IX6m�O<c��C�OT0oZ�6ȡ���Ӵ��5.�$�V�s�4V?R�4�;R�J����<QU��G��ݔIɴ��7O�I�ʔ��8���0DreI��'UF���w���*S$�O`�d�O����H�˧Y��C&�F47�8���Rr��`�7�C�T�0a��?A���r#OX:��M��]��dl�2�;j�(�@FC�>w���ٴ]R���ڪ�~2��Ll��OF��3�ϝA��B�46l���D�I��ԡ��C�y�a�6lRA�	D�m�/O&����H�(�Q�����w��cF�;LN��$,�����䟬��dy�C�?e����'���'��I�͏.l4��:4��>6ּM���'�J���O�h�'�L6�������a���Q�K
ZR���0`K;?v�X�Z�S�n���<O�(Jp��:q�nq)�.�!�"�'�B)kd��{�ӡ���2��c-�LJ�������I'd�h��k�̟��I���Ԥ��C0h]���Hp������Aݟ�Z��l�^,�'�7M�O
�hҔ��]#7fZ׍��fH�(�� ��LP45���*��q�4'�Z9�`�'co��C��<A�@�.�{k��#%,��gP�L"�1���uF��3�lXy2��Oj$���[.`���Ov�������ģ��9��kW]kO0��ˏ��RapLc�"�?	��?q�'X(8��+ON5�愀�*�X��DE<\��*��EB}�BbӔ�o�<W!��I�Ȥsқ?�Q���}kHEkf'֑r
"�R�j�>t3�Y�''��Q��	+ں
?�&�|)���Ҧ´$� �DC	+�.)�DH�,6�G�̘T6b�'�2�'��Q��sp�Pv��	�,�"�CsL�dk������o��I�MC��?%��'���_$���{�f`�p,��u��ջ�A�>RXUn��J�H2h��j�rW:O| :�Ҳ�ub�˵TS>�{��xzȩx�˒�Ff�A��cQ^x���/ w�>��?���
�&�>�����g�jh
���(�8��-rcn��<���?فɌ
^�"��'W7��O��>O�X���GIÚ�5�'p��x֋�b�|�I%�XDk��̦瓓��z�O&#0�r��T��o�!A��(�Ê ?�p�oL59�B�Ԉ5L��N�����"L�'��'n"9"�珟�>5" �#'�,�4�'J^��Q�ESr�x�������?�b��'���p�@f���!��b[�F��	0�M[մi�6�:�(�O� i�^���� F�'��If��)�Ņ/U��aQ�G�C�E���C��B4O�ԫQ�?)%�Оg�剐����i�(�1Pg��#�\���&E�R:�?���|����?�)O�0R0A��2�Z��#_��p�c��'g ���b����ش�?iǋJl~��>i��i��� F>&���
D�0wʅQ(~� �p$G�6���v$V�$��9s��Yw���8co]�<IBO��7� 1�um�{W`Eb�����$K��n�r��7D��?����?�'b�j)�,����sOa�|�X�]&�.�S7���.u`�6O����O��ɀ�_���'�M�;`�
���?I����A"Y�z�!2�i��6-S�b~����,�0�ѕ�?�:� ,{�U(�+�
yy�Սq���r��1�#}�$u��O8����|yb��O�(Q���,f9��X8J�a���]S�X��B�w?6���O���O�l]"�Ó�J�<I��?q��^1k���NFxr�0��ۏ�?i�gG~�
�>i��i�7퐞}!\%�	4G��SM9{�@%�Jx9%��I�9|L�T��B��c�Z>��se�ON�@���Jʦi@rfH6U
�W��*��x0��?��4NH�1#�U���'�?����?�2-�z�V],$���^P d���^�$���EP~B�z�r��O��i��4�I�]v�iS�b��u���0F�p ��o��M0A�{����ti�x������(eb|�Y��@�s䴬�V�]I�]J��[ka1\�<��u�Nl: �[�?����?�����I���E$- ��v\Z������ę�ne��1O��O
����m��ɔ�\u���(.�X�k'�]>WRl˨O�am��M��j�m�/7^���O,F�xŌT�/:L�V5
њ�Ek<�J)�fD�:�y�MO!$�n��I:%F��/On��Ʌ7�2�O^���Q*�FBEP��3��Iޟ���џ��Hyү@�[l���'�ؚ��8p{,��C�)aX� �'�H7-�O�hp星� �O�ylZ8�M�0�N,c�\��V��ͮ�ȓL57��p�EƐ�ҿ&%��LN" �Yw�֕��l2�V�v�U�ʇ��%�&+D�:���'�*x=H6!���՟�Se�}'?��_�x5����Sr���`X�q��ß���*o�^�!� 4���i�b�N7�y�a�;K&f��фǆ"�|�x���1����'�:���7��Ok��#������ٜ'�������gBS��5rAE�8Sex�ϓ=W,m,O���I�sY)�o���I՟L[���]�x�P͊L����p��។�	SyRf��5��Z؟(��ȟ���1,L����� ��C�a·��<¥�)?�V���	䦍@Q���0Zf��#������1|����N���q ϖ
;�����gǿ�F�Y���+@1�o�
�oe�x��N\yթ	3���	ɒ#� ��7d��5�>�D����څ��O��4�:��ON�p��<i�P�A>ȍ�"Y�M#� {T��.vW�:���?�p�i������D�Hyr�i� �`RE��u�!�s&V����u,b����(�{;~xQkA9p���d�	A��cXw^���L�<q���(�ڣ�R��06�ȟL��ޔ��� ��?����?�'� x�,�hL����>��@�%<�Dh@ ϯKR� H#��<Y����D#M[���k��.����c*m�ڔZ�X����ۦ��4L��=�o�����?�d�L<Nt�J�(y���	�c�)�N �*�qrt����-,F�)U���'���$��l�VYZ�&�O��;L�8\�@�Ѩ,w
�UN�O���O~�$�<i��A�u3x�ϓ�?Y�`�l�w�^�1�*4@�̉�^� �����'����?Aߴ�x]���'��!�mE
S����ɳ����c�6*�R�ΓI8f9˖�]=��S��m�#S�?wH�1G\����I�=	��qQ��.kf�٢��O��O��i��̊ej�������O����P6,B���	���g��Ae���ʩp@�+��Tڴ�?qA�m~�w�^|(�aC�?0΍u�_�!*Z"h�4��\Xc|���'�T�����X�x͓z��`Cnuݽ�q��0J���+c�3cf�EFQ *[Z�"�W�dR�b���`E"X;�?����?9��uø�z���w�N��RO��Q���8��Y��B6'�0�P��O��d�O����TN˓x������Ǒ�f�c���~nl���[��y�4FH�����~�/��6P���O�B���Y�3�0��`Zu�pq;@�Y����p�Ү�y��Ī|���I>�ؤH,O��I�,8-{�ƚx0a��ۅx�QX��_;o�����ڟ���̟,��Ry�gC�<��`�'��aP+��*w���YE�5j�'G7M�O�� ���<�OԠlZ�MKV��d[�#��1:�m۳OZ�m5,2S/J	��CP�<��
�"G^�]�V��1�R>�q���D��	Z�c�!` B�!_�(�c#.I�)���OJ�d�O
�)��^߀����P
/�<�5@L�[b�����|���O����:'��⑟�k�4�?i�'�<A��D��N� LTq��)��A輨I��'�Db2�Ƀ:��O�4)+�$�(� �'�h�"i����YW��Nze����w��h�ɕo�&�-O"P�I �JЂ&�Xݟ����X�����R�"��ɊT���a���<��|yZN|@��CM��?����?q�'-6(�0���t�� ӏ�( ��@�@_~�.�>A �it 6�] y��U�:�و�O�6�+�+Z�a��v�q3k	T4-r3�@#��)2��B{!����](��'�@ԥ�<)��q��t A/T����
1R�[�.@���'��On"�'��	�x Ð�_�=�R����[4+Xd8@�)�s����'U�6��O2�q��t��O2�m=��kRKҖ~�Ȑ��%�z��۴`OZJ���B1ȕ0#Q�<9�K� <�@��~��i�P1OR����D�.� ���;
R �q�'vD�ՠq�ѡ��O����OX�)��P��ʧN6�C�Y�f`���ڀ��f���>����?������Đ���]�B��ReV� ��� �Mȵ)��t0�4I��m���~bl�-,��Ox��PbKJ�J6<��-Y�P�T��ޚ-�,eP�Y1�y�+W"o���	0�i -OBt�	9,p��k��� xV/�L�|��ƍ� ��j&��ҟ������	}y�֥FWl[�'�r�'�2�4�q�Vu��CI0`7Pa�'���O~��'1�7m��@RE��`�� ���W�%�����/4`-�磘�Mt�D��r)�)Q�D�t�
x�_>]Ö��O�!��%�=H�͕zҮH�',��XR)����?Q��S��5��ϝ����?)��?Qpȑ�{3p�#.@�c���?�5,�,7[���(On��\H%�!?ͻ	�d��6�E�c���� c�.D-����J�3��Q8ѹid�I����p��(�æ�y!	$�\h��u+|���׎=\��c��$�K�C�>.��>]�ϕ]�����''��'���J�51��U����"��;#�����p�Y�!�� ����矰�	�?�
��I~y2�:H���T=';���{k��x����o�I���O�C栁������:���*X6njh�jc��	zboQ�]t��a�?O< �ܪ�?Eo�#O�剻�?�D&�-��51��ѳp����q��,1g�0nR �?����?���?�-O^�U���0;�����bh;জ.�n��% �V������	7&�D���	ҟPl9\f����,ɯ0n����m�x�[rRi+h;!�Z�X)��I�. "q�C��Ll�a��������1�'X8i>]�ɟ G�Z���(¯U&�r/�ʟX�Iş���Y5P%?��9y��툄�H�|�Z�g��,Z��IΟ����#�4�A��!"G�i��	�yB���b���1��8l�l��RBR':|��'��3�h�b���Oi�%����B`�Н'!��*�Ƀ%<�A��-ӌ�~!��	ֳ<�>HΓU��-".O�	�QjeF����TӦf�D�0�� Y�R�x� T�����Vy���.���p�'Z��'-����7A$1)rǢPr��e�+3����O��'s�7-����q著t�v��)�)�/:MrA{c݃+Bܨ�JH�<����E�&�90�G�UT��O�H	��v�Lq@Y�4!@'�4,&����F,v�9e(���?�B�h�m���?�'�?����	�b��}���Wo�N�y��:?_H�1��
tt���'�v��O��'��f��!CL�5���΍���P#�6�I2<��ق�CT,t�,[R7O�|S��Z6�u�ˉw�h�1��"��+;��))g#��L�Y���?��c�-r��hr��?�����/ڟ��W�f�*��7�6i���`֠R�c�dX'E��Ot����p�Ɛ��8����"ܹ-���a�.x^��sa�@�)��gcӪa0��ן�-�C��Ӑl�D�1~0H�Fj��t��Ə�o��z�(}�l2b���i��/\�b˓�ҍ�"&�"�6�'��	R"
/q��KqFD�f2�q��'���'&�U������\�h��֟�ɍK�^=�ʆA��M�T�_���	�]���c��	��M�c�i4�rvl�O��h��?Mh3��U%dS��qՎ��yќ' ġI&��:=Ra�d�	���醀��Ê�I�<��sH0S6�^N
�k����	��DjĮ:
6�'?������	 �a���6%hE��|��&.�O^ �Fk���	*�MC�U����y��El��O:K0\t�F�Nj�<�0�'ܓ:�6m� ��-`�P D�ڍ��6Od��gOĜ�uh�*�" ٺS �xya�ߵT���A��vy*�O&m-F�*ވ�d�O������� �1Zn�a��T�>uqB+�0K�����\��BVv~��'a�T,�����E�bH�U�.ݍX�fq ��A��HՕ'3��ia�C��O��1�)�#����6��P�V���H7�A�_~�L
�����l�@�0O�ť�?��ּk��ɟ�?ť��s����8eVa�7MО-]ցp�у�?a���?9���?*O���ŢԪ3��d�Zw��{�����)S�/��$����I�Y�4��I��M��i�Z\�0'��V�������C���<S������2F�'��98U��Ϻs��Ϛ0��˧,u@�>5(B8p�� �6��!DCߗg�𡊥��&�d����x���?9�U��x�sޑjEJ�I��0��L:D�Q(h���Iݟ��5�ޙ<� �z���'��PI�'��嬂;$Έ���$���1���,�(����'�z�k�Lh��i�O.����Al��dA3?�� �]��r#ʅ���C�'H���I#)0 ��(O�Q�I� �JĐ��^���I՟�ѡ��y�,�`ɡ(o�$�Q��?�/O
<���[���� ��0HT}���){t�C#/�d�p���a;?i�V� �ش;�֊�*UM�����u'fd>M;RIЇh� t8�O�YK��
�(�60hc�G�ڶa���~��� Tu��	&V��A�$���M�'4d 	��+� VUV]i�'\l\�C������T�'d�_����R�^u�	A�K2DRh�,���'?9Ҵih�m����YR}��m�T�#�����݁��'��ԁ�IE���cŇә{\ұB�$ v>��92�:��õ�7M��yBe@�
	!KڑzP�:6g�%�?�C�'_��qEOݘ��E	���K'9D\mC���5d��o�!*9��uP���	�?��� -����y��ğ]�����db��',�H6֦͟ͻ�̳��iS휋P���D@k	<P��ؑ���J�`Dkl�@�bK��y��)t\�y�Idg�� *O.`�ɇ^���I��p�<��DšC&�� Ԩ?
���f+O�](�ቁg�B��?�Q�<�& �Vf�&20��Zrn��?Is�@~2l�>IP�i��6�s��J�"��X�J<;P�C�o�>v�(1[3�V�y���TL�E�R�2��f�t%ʽ�?af#ߍ-4��j2Ǒ�C��Jeē""��ߘ'���(��<�0<��+,w� x�̉�+�j�ʷL�<�?	UjC .�V�*O2�n���bׂ9?ͻ/��Bт�V�&�ӄ�0����"oϻ[� �kf�ir���I�s,`)�����yr���;xR!����I��:���c�R�1TL��i i�H�B)O8A�I�^FQ�&�>�i>Q�Tl�r4�m����0XF�Psh�g���G\�C&���D�O��I��-���z ����)P.m�fƋ#t|�0��O��n�.�Mk�n�h?��K�8�Z�'M�8�NB�NnfQc��A܊�!��v�.��a��<),��,�t�D�;mpH�'i��$҃~��2bM�}b}Ѐ�)UA���C���CCaz�Dљ'v)��'d\lc#�ȅo��Z(c���y2dh�0�d�0,?�ɲ���O:6��['� ,��#Ø��X�t��,5�zgN�+j4�l��2\�����^w�fay�E�v��A��(`�«욭Z��ɽ� �{E�ʯ{"�jV�4�"���I	/oq��R�Ph(8���L�w���'�r�üY��-�ȟB�n�����ëy����mđA�*���/V��#.W�|���ɤe;6e��a_ߦ�S:]��#���|p�I�H�DQaiP�9Y���섒�h,�0hW��;(N�"Y���>�8�t�'�B�'l�5�4��i�	F	��B0Xr�'�"Q�8�UEL1XU|��Işt�I�?Q���$[7���w�W�:�d���J�)(��*q��ԟ�nڸym������J���@jXV!�5	˴P"�� t�^�U�A��K��J�X;�O�y������4~���x+O��*4&��S�B�`�a+Sh�Ce�����+��>D�1���������	ey/U9&l�����\g�.izU��c8-J�]1B]�	��M��q��'���A�����C�L�R�ضKT^]+&Eʅ	H7��~�&I�c��8�h�9Oa���ug��Qqp���pՀ�l˯z����"��
4	��2�?�4�7)�\����?�����sN���WV�%����Q��}!d�T�-*��v޼�$�OZ�d����b�1����[��]"@H������ {�v9�v`Є�6$�4���^��~���I���OM(1	��F:#D��@/�"8��/@�ͻT� gT詝'꨸��_��`�ة���X�@�ER�i��i�ɹ8��H�S�=v�cDG�Ov��	ޟ0�	���'4�D"� Q�R�'����1i�۴f	}_N\*�%.]�Ҡ�yB�'!��6D��@iӮ�x&�O� �a�p�>������|5.���r;�	��'�v��w�+UK�y��,����@2��%��E�8�uH�Q������\�=�Az��۟�I��8X"�.`9d$?-�	���w��tbc�ڟ~F�h إ@�d���5 w8��wϟt���M��D�����?ͻ$T�MP�/�o:�Z�@G�>FȁJri�j����ixp ;~2�Ls�"�:�y�`��c���;*��8{hڻX���#��E�b��Q!I��˓(�ۭ`��	�Q�'��'����U�\X�Y�B��>_�MGk#s�����Q�L��F��A7&��	ǟ��I�?���t>Y�	t4�@� Χ*���4$Ǜ;��`�O>�l��McS��|?y#�M��!U��'n�%d��a��Ƀ�_��E~�a4�m�@�\\ 1+@$�O�)�TK�ry2#�O���>8�HP�䇣Ę���(��B�Þ~��$�O����Oj�ĩ<A�	�?1W���wK<���/�5I]�L$��/.�!��!��F�'����'��c�>Q�i�^6�]�=�T�@K���V����K�y�����D��5�"� �ѤPh�pXw�ܛ��`��*��q��c�v�!�a
F/D^��s�dę)�У��O����O�iĐ)�t����ǟ�� ���t�����Y�)�t�$�O<�Ą'bY��8����ꦹ���/�$��L��4�WmǦ.TT����	ZV��D�����' 6Z,lz>a�r�L9.T�ER��~��10�K�4�d��hѳb�E-=j�IBS8O��3n�<YA�'.�`Sv�Er�'��@T:o[P3�@;�^�����9#K��'J��)}�`P�j� �I��x��66�	
���'dD.8	f��
Y
#M+?1V\�X�4!��FIY:kƈ�dP*Z���{�O7&����;u�Eq�P�{�����Ŵ�A� �?� a(��RVȋܟD�g����ƻCp�i)PM[?cՆ�2u�}�<a�I�	�*)��<�i>9�I��`�'�V-��	JD"�*BI0n�SA�:� \ �Ob�l�ğ�ɥl??�qS�$��47ֶT2��'/���rd�Q*�pT�iKB� �E�/H:աP�S��y"D[�r�5�;NVԭ�G�d�Lq��x��&F�3�&=�e��O69����|��g���@��͟��S/f�R0�OA���WE��9�'-��h����݊�F8!�'���'H��G�'�����*D��¶@A9u����0H��;��-c�4sܛ��z7>�D
f/愛ʟ���w�p��arc��i �8�5�+P���!	g(��2!�^�b� ��`�R��H�t�F�C E��?Y�cԲ��X"�'�M��7!R|�B�'���'E�	A�<�A�&r������9�! {��ݰ�!�A;Ll`�$�؟̠�+"?��V�L�ڴ���!#g����[���l��bȖr�=���$��d��'�y�g�,e����@�Nf q+�ĕ�C�'����Я
yꮈ�0AX&GV$$3P�x�" ��韄�	�|�@a�@]�����i��"'j�DS�ِ�C8�<�Bn��T)�È�R�����F�'�Й�O�.@#\��T��A��XD�G�O��s7��P�شl�����;�L� >Fs�i�,�b&��O<|Eq�G�9t�,A�\	NBx"�Y ���!�9X���� �� l^�E� ��/
H#4�Yf�b'^�X<�q��';�����ύ%&iB�Y�$�`��˂o���R�W�K���L�6�p���*8R6�u�l��=�F�C�	�\�2/^R*����^�o�"Lc�aH�&�ʕ��$��'��EYF��?-��ˣ/[zz8�#�Y�s�4���k�Cf@�R�}��
��\�d��_h��	 w����O^�n�V��d��x���⟡TӼ��G�̒(c�j�M��F�����=�"�8�A�7+�1;�@*J�6�'&2�'���f�<Y�I�0I6���HO�G)@a�N�u(�	��ڟ��`�,�'mɧ�)P$F�6�w&��^��7���K%^���O(���O����<����|�`��0T�����`]6ypv�9��o��Gx����'@�ee�M��=��ʑ?�Fy��D�Of�$  |����O���7���D��K�����x#�i�T�YN�ࠛbe@+�"<�r��d�'���'��=cbܻ�L�3�eS��8�	d�h���i�����O*m�q=��D�?Q���O�����N�Jc���M��&�*�A�&�$D���	���IΟ��I՟�c��ޛ��@���P{d����f��'\v4���'Q���~�'�?��'!ظСJl|�q�H��N�D�&�iŪ�#�O���O���O���M
\���(7E�I�`�Ю]�}���W R,V6-�%}�h�D�O܉#��O�T�'k��OӨ}��42r@�� `��=v�Y	��j��'�2�'RB�'��)���S쟌� r�:��\��\���׾�(���iF��#�~"�ۣ�?9��zumA�ɷƔm;��D�j�pa��A4q��4�?�����$�(\$'>-�I�?YS��U�$9&�͹Nd �`t��W����]���D�On���(O���-��,ec���ez�t2�i�剾#�P���4�?9��?���z���8Q�<�@���T��c�G*$�pP���l��(u�"<��F[C�ɶ$������}��Dq�dB�k6�(F��m�<��ڟ ��	��D� �$�"0O�@��Կ-uz���<Uqm<#ID��	G�IR�c>���Rz�$����<O���ڴ�?A���?!6Y�yQ�I�`��Iџ@;#�gӦA:0�H&� �P������D�K�1O����O�����> ��+���(9SQ�vҐ�l�ǟ��������ZZ�$�O��Zs�O�\c8"����pd%ᶀ�
oJ��']tu ��|�'d��'���&l?2�Z�� �Y���p�������K����G!X���O� *q�O�4�'���H*|6��v�*	qU&��t��hr��|R�'���'��	�EF@��OV��c��D��$c]����ش�N���?�%�A�<a�'�?9�K^X;�Op�X�hE���cU��
�ĒcP���	��\��\y�)�~D,맻?��(ڐ�ۗ�74����d�����'��Aq�'��B��?ѷNP���'ڡ!ď��^U�4!��`,����ןH�	Cy�NL��'�?��BB�;Ny2�gD�lX K�[����؊������.MC��Z��ΐ�Y#+&O��HbN 9L�luJS�i�剰Jm����4�?����?���W��ɬ�l\��7�<I$���"x�e(�ş<�ɝ)}P�?a��QD��A1�pf��;Le�{���Xg7�>%Y�Qo�˟l��ٟ�S����[�Bl��|�$-���U0�j�*tCI/*A�qm�J�T#<���n̓�?If��z�B���ᓇy������p>�6�'X"�'���ɔ��>���<1�w
�n�*�V�7��$j��i�E�E.O�Nb�<KA�Ps�	�`�����[q�/.����D��v����q�iAٴ�?��`O�K���!l*�	��Њ������<�(����d33�D� �f���V�T��Y�I�(��ޟ �'�ȱ��癐J̆��Q,�?��T��)]���`j@���?�T�^j?��䟔�	�~�9$o>~w�]9E��ª�ȴ��џh�'3��'[�U� ��'Z7��d��_z�t�W��M)
R���9�?!�lן��ɠc&���|�/����ٯN�� �EEQa�6:�<ђA�'�r�''�\��I�m���'5 l�Ad��-A��UR���q2��i�h�#�~2���4��$�O�/n�P�JF��'Zw.y*�.�< 6-�O��Į<��g�1��O�"��56a���nD� T9K� �@�(��,�ɢV��˓;���Ox��?�i݅�O޲l"`�yd���y�m�>�^(��k���?Y���?1�'��$ H'��i�D�b��x����;X��
��OV�6{��Ex�)�)Pw��pa�]����&̓V�fi�lB�'�B�'���V�T+�gb>�����`���)�j�((�|� H�?ɡ � Rx#<E�$#G�5@�p�u�����0�V�N�A@7�O[mZ�,��Pyr��&���8O��I�4il"�ueR�}^�YQmǗCf*Xh1ቺ��Og��OH���]����K^�y�.M��i��ʴ
��	�7��<�š����C0�-�,ҹbY�s��uD�!'����0?A��?�����ҢS������Ҧm�̱�O��"Up���*�Zyr��?��Y���O��i�9J%�0fo��c`��Gd2��rӸ�D�<1��?�����d�5[;�X�'t>�Őd�B
2����#�><c(����1.���O��I��O�dQ���8�!�Ĝ>'�`@���#/� W@�9����O��D�O�˓x���QB������VIq��&�]����[d�7��O�����O�e�PV�����~��Ҫ1�F�H���O��ث����������'r�X��5�)�O�������_�j��!Ǭ�7QR<�r���<�f��������?��yZw8@���۹J}�Ca�Ά|���O��$��kYP���OH���Ob�)�<�a$�t�`���,�6HǮ+�L��;�Ј@��yB�44zEFxJ|��DQ+:��L}�aôHY˦e3�Kղ�M����?Y���aS��#�<��I#�G�;��ը��Ղ6�����
Ŧ�����IP�)��?٣eӫk��4�I/W�t�QGI�6�f�'���'12y�E�>��m��<���C>�EmZz!z4�eɜ]:�	E�[��7��O�ʓ{%�1�S�D�'�2�' z0��׍EƬ׏ܐfI>4�@�~�p�DU�J�
�ק���z�,���e�P�I�?�X�Yz�SQ� 4/��T��r"��@㞌��ٟt�	uy��y�u� &�j ���ȴ9��
��d'>��O�00W6O��)�O��T?w�PMf��{�T�B@�9IJ@���D�O��d�O�˓3��@B:��Xx�HY�J� (akM&��ٱ��id:���'D�œ��yR�O�R�'�l��OrYH���]#�jԹj��*�i���';B�'$�	�8��s��X���1�J�>pz\�ꥏA�4U}n����[�Ez�4��k���I�>��|nڻ�\B!�ؠh���/{xr�;òi�b�'��I�Q�Ȫ�����O|�ɟ�_躹!�Ś)�N8���ݤ�}5OXXx���O��I����OH�r�n�^�r���0s:���Z���[�TB�n�7�M����?	��2Y���	� N<�b��k��}K�V�;���1�<�?���5;����?�*O�D����Ԥ���0��aAQ�$���M��U
����'A�'w��L�>I�Ņ�<���փ(�B�Q�B�d�hB4O�&n���n���y�|"��8��O�r�J$V�d�:`�5fyi ŌW�`7��O���O�$�o�l}b����y��' r*ܴn�� ��& 5+]�e�A��%�.Il�^�IUm��)2���?����Msu��.,3f@�־u[���`�L�$r��'F����'��/�yr��56O�Lt�f
](�)�J������O���O����O�4�y�`���#]����C�X��(],v��	�6�<�	��K4�}�D����ɒx�V�����\�	k�C��9]Љ;�ll�ؗ'��'n�O�
���p>��Q�	1`����>8P���dn��XS�5O\�d�-����8���O��� Z�xx�N�g�>�3GJĪq���v�m����O����O��~Tv-aR?5�I:9����[�"5a��1;o�E�ߴ�?Ѱg��<1��Q(�?��0���'����q.IB��[5=	X�8BۓMN��'��W���7�;��i�O��D��(�ӫS�4��Aȣ(�����r��b?�"s����O2�r;O�˓�?�G3�T#��]�D�L��M�>�H`#��ie�I�K��Sߴ�?i��?q����I����$��< ��1�4�G�j8�T������� ��Iԟ��'�u�I|�w!�`�� �5�Z9�8H���ۦ92�kP��M��?a����P�pX��a�䘲��(s���Z�[��A��M��<a����F��1���$L�$��1`2O��>���6�%n�����ǟa����D���D�Oʘ��iSH<���@�8u"��Sb¬U�T���4�?a/On`ڐ3O��㟈�I��8�@��&7��8B䍄�G�<H���A��M��(�p3�X�4���q�$�I%&��	�?�؁I���s*�  �=*d��%;�(�@��e͓���O��d�O�˓lH�a#!E÷(6��bA�+/�p�q�)V&nQ��/Z����<��+{�L��ן8�I�.������ܩ��zA,�E+T��e�5�П���ş��'C�a{��w>ŝ�g*4Hs,׌Ki����vӶ )0OB�DO���D�V��O����Q���B�p�,���&N(���`�^�$�O8���OXʓ�z%��X?����XYw�բ.�r��tV�޴�?��+�<	ぜ�?��I^����D�8G�lX�6g�5Yx`�P�ʂV�Qoޟ��IOy�mК{ު�'�?���2a�K[Ȳ�%/��%��p�R`Y�
JQ�Q<�eS��?��QY~�T����w{^t0ǥPD��G��.����4��dPb}m�ɟP�	˟d�S�������$�vF�z%fY�2�
>�z�����O����9S��O���O`�膕��j*���"̻�L;aŚ��M�q��a{�&�'�r�')���>1�)�<A��ˊjz�P(��R��-��)v���G0�y��'T�5R��c>��	!R�t-��	�T$���ShP�_;@!Zߴ�?i��?Y1�:8��	�O��D�O¨·i���ʱV,�􈊒q�A�ߴ����i�`���'o��'�r0��D/���i�	.U&�T6
}�|��ńJ�̕'9� ��?�#B]B�\cZ�u�FG��M14�#�
eԼP�OF�V8O\��?���?y)O�dR�K'D 2�L	_8H�+D'��������?���LVx��O �'�|�XEH��*���E�gc�U��LJ8�y�R���	�4�IKy�B��b&��Rȉ5�g�ᓅ�ğW~>��R:B�b�'�:�'�t�'�����"E�=�T����� *�`\ �R<]���ΟH��ʟ�'O�uū<�IO7#���j�E��
B��-A��n�ퟌ �n�� �1A�On��)
���d%}�oܕz�z��`ިv���j����M���?-OT�ҷ�}����ӑz��:�&�%"0�Ĺ��9�N��Iw�����Ol%�U��,�y�dY0V�h����۰m����� ��M.O�mz$%Aউ��������	�'Y��.9�H̉ �ЖVۄ�[D#ѥ�?���j� �`�AY �ħS����DE˯g�~<�"j��{��o��=\��ݴ�?Q��?)�'��IDF�q��a�)��x�!��)RF�oڡB����u�����Ol��&��j��I8͚	_,�H!d��������\�I-�RA (Ob-�'��Զ�M�%r��a��E�O�D׎W��]$�̣�Et��?!���?�p	�F��I��a�I��Fٴ;h���'�� x�M�<��	r�X��2	T���C��T�QL�pqrcS�bچ���	}�����b\����۟���qy҈
,�>�'�VxxT�0	�|����<��i������GW���?����\ܡR��$r>h�aaA��x��q�dH��?/O����O�$�<��@CK�I��YV\�BcOо'ڥJ�0� ��?q�U����b���?�@."��d%D/�6�``��d�њ�i2	��D�	�t�'�s��,�I�:w�+�-��t�qY������n���N�P�r�'Eh�ə'\�wb(y�o� �
h#��o��o��	Ayb	��|������yـ�ŦEOf�!6iيHY찧�ۃ}m��N�'���'�bX1�'��'����%=���EӬ�4��D
=<�7��<��%ٙV&�怼~�����RR�yd�P�v�b�S�$��|���N���O@��?O.�O�x���$�~R ыR�)1�%0%��M#%ʝ�R���'��'�t,�<�"�w���Ge��$����"�t�@��ǂ�M�Tj���?qK>q�K?�ß��΁M�(8�@ռ���"`����MC���?���dh\�`\��C6OP�d��*��� �ذ7�)��p"!�[�)`2�i��'�Y���)�O�$�O���bL�N�!s�.��W ��eXӦ��	?o�d*)O&��O}�P��i��A��*I@@x��ٸ���L<������O���ON˓`Ѭ��j�1��H{�;<�0��K���
)����|���#�?�y2SO��<|a���מt#����!Jڦ!�������՟�����ؗ'،���Km>��W�P9^m�� 5!h�2 `�O����'�d�~��<�(�V���S5D����,����������'�2�'��W����l����'o��b 獐V-��Z�bb6�P�iM�d��~���<a*�T��3}M��)?��!�ܕ9�f��0���M���?�*O�\�UGT���'d��Oڦp i\*p� �=9�Zт����yR`��< ��'�Bq�'"P�Hq�w�~$Q&hY+ᢘc#���V	�Q�4��$�~�.�n�ݟ �	ٟ��ӻ��I�B�`�^e:�]��+D˔)`qB^��?���k�����hZ��'>-�,9	<.�����8^�m���c�(��4H���I՟8�I�?I��O��2'7O���0M�j�"�a��O����'������.?�*O�|�"���O�|I�+RpɸbMD�y�x��ަ!��쟌���L�Ty٫Op�870O����0^v��ٳ'V��-J�&�r�а`�/��'��"�y�'�"�'��H ��2�F��ᨈ0�ޠ#�Gk���ě����'tH���'�R�Q��yR��5V�G�@h0q�"4"�z��B+��M���&J̓�?	���?��?)O`�{�@(Ͼ�9ҊP
'���3$F�
^���'����'����4�y��O�"�'7:��B��6�x��H��	�A(��'2��'��Q�T3g�R���DN��P\���3������M����<��^�<���"��?�``�V}" ���E�'ѷ$?�t��$ڷ�Ms��?������O��8��|���/#�l�<D��M��"�[6�O"ɳ7�O�@��'���OJT�hH<B�\'9K�L��{��k��7��Oz�d�<��A���O�b�O�:Ygj��OBV�B� �$Oi����%�~Rƀ�?A�'��3�N���.�d+*��qiA9�Dil�[y�����6��F�4�'��#�<1���o��}y���M����b��.�2L���<Ղ0lO@ȶ�۠,� Q9F�PW����id�E��Iz��$�O����D�'���
��r��jE���z5�U��, �-W
r�i�0���ĕ3�1O��䐳DZ��T�9O�|�:Q�@
9n���k��D���E����'n�� ۴/?ڴ�G�'7����#">����>	$�e̓�?���?a�
D�I��L�P�>��!4N�&[n�&�'`�PH�>��A�<��K<���1)��Y�7_�%~}k@C�JL��'R�D�ON���O��D�O&˓��E��c��W��yS��W�d��@S�� 8�I�MК��ҟLI�`����(�ɝ,����\t���Ŏ�Y��Lps�,�ğ���ʟ|�'j�9��m>��o��F���k얾]�p91��n��a��0O@����9��$��F�$�OR%�pX�ᶭ�1V����1el�a�<���)ʧ+0��;f���q*:ԉ��êL�J���+�vy�!�����]�㫖�]�e�?�0��/
[�P�2V�JF���0�g暠��)u�����	G�,��	$��<W���A'�R���4j2IR�v^|��l�J�ԕClA���%ȧ��"c�.8 ��_�'�NT��LY^�<�V`ՒL��%Hri�#6}X5��d
$I� �HS�����!�@�
'7Z�Ӆ�AM��I��X���SXR��GA�${� 
�2yE�ɺw��"�4��[9p�2����?Q�N�$B ,��?i�VF��%  u���"�)��&ζ%(�mS�wf@�xdj�6%����'r�,8��U��ԝ`FC���h%��[	��'T�)��,���0^��P��&T����h���/�!�D�<���q��<^P�I��'6��,S�#<���<!eǋ8]�(�V�������+���?Y��L��q�1�[��?a��?I��H~���5��?�?a`��c=t��%>3B�<#s#l?iSeF�g�% FP�,��x�)@F`f��coǂa�Vp�n��~2�ۃOTʌ�ԄG@5����8g�v`8�H�!c�'p�X�4n��| ��OR�D4���d�=%��hP#�g��4ꥍE4/�a�{��'
��A�� ��S��X�T� M�#<���<�(O�9B�hϘ2Ƹ$���8^(�����7Wtl�p��O��D�Ol��˞*���9ף�Od�ӣ;#J��aƛiR Y�3�^q{��O�AG����(���=I�n�(�Ry�Í'N#�r�,Լ`�#Wk�\����'�'�l�A���?)w�4L#�\ �^�S����eK��hO��?���9��	c�F�p� 5�0�Y�'d#~�'�X��x[1	U�[�('	�<q�C��<��}R��:����+�;�-E��&C�I�C�ȑ�ëJ��=`��-bBB�	�GJ<�:IG<�\|kE̹6*�C�|�@J�lĲnx6\`1�ޅ~��C�	Z8�L���D0P�c�z�B�	{�ZuM-����%A(EcnB�)� Ҭ����v����!��1k�"O�)�e/���X�fڛzN~e�f"OrȐg�
5r� T��D�	33���5"Otm�̻&�J�z�n�H�򅹧"OBP�c]�IB�sb�Gr��iF"O� ��!؀Əz��й"O�DKA�/��h��mݼ�@���"O�\0F� �JRٺw�V05�0�"Oꈻa!�w�4�boԣ{��R'"O0Й0��ik�u�R�\�O����a"O����Q^���&$�+�NI�"O�H�� �wlN�
�c܉^��Y"Oซ��E�ol�a���>w�yYA"O�yi`̃�t�ĳ¢֭L�.xW"O��E#�y��]��Nүp� �Z"O�Ȫ�	��ps��Zp-�5�`��"O�Y�eN�@sTU�Ы\�q���K�"O<QxV	������K�JD��;�"O�3S/ۓPJ~T��d�5@N\�"O��CNF�HZp���"��fL|i�e"O�<2"F�\���p�E�/1��C�"O*hip�,0j���%Ģ�+g"O�|�v'�*G�T�x�*҉j�dB�"O��(�!U�e�0)D�g6��"O<�3	��h�rT�&��?x�Ȧ"O��`���4V~���G�4}̄�&"O2E��$$�����&�G�nh@v"O^�A7e�v�t����C����"OҨq�ԵWϺ`1�$�|�T� "OL(iw!�m��{�F�� o��"�"O�(�1, g���gƑ V�0�s0"O`$8'���m�ȊG&ކi��Q�"O�!x�"�,	���ł�n`�K�"O�Q�R��yD��p���(V�D*G"O
E�uA�wjb�c@͕pW��h�"Ov|ځ��IM�}'m�o, D�$"Oꭻ�΋�q�e���� ��Q"Ol�&�Ow�!5������V"Or��w��(9�]1��J.���"O��bf�U5L����3g�*L���hu"O���5EҺyjHl�S�ݾi$�I�"O��3D�K�������[瀽���'�~�C.O@�r�m[�_<
ec�	Q)P(��r�"O ���Aϑ6I���o������ɸkq0�D��
Z�g���C�]~�2u�B�]�yRџ�ീ�lX>y�f0k���9Y� �yq?�)��@����Q."���*ބ �/D�@���1A+4��+���$����(��X���@��E=�-ٸ�]�UO1�O. S�M�>	��U��;�c�*�h�ѡ�`�<�૙�y�j`�M#�A��
Z�'����`���M�a�)I�y�
��Z2ybB䉡5��(V� =�� �Yq%X6�׃��"~n�?4�\��gV18}�8����00B�<=�D���C�M(�d��I��8%B�	
��i
B���ڝ����160*C�	?OS��hĬ�E ���Ƒ�"��B�I��"�XƬM�|=��s����L����I���'�8��M�5���f�_�&�����'n�Yz���Z��P�G�;3O�uHK<���*�S�'J��Dr��8_G�4 ��I:R\����{����	#@J@���n�x���<��f�:8Bay�+ӣ@0�T`�	?�Qؕ���x�#Ã ����% �ފ��D�
	^Ȅ8�I�O(<� �u9C�Ξ"�����.^������'��{`��]ܓ}��U�4���5\Z0	�*�t�"OH�I�˚N�ɗD�3e�ܸ@�x�'��'Jc�b?IY�d9�%�4� `p��S�;D�0,�*��q'��F>��a��!������ �:�>�O�`BDѭ$�Θ+0 B�hjJt�ȓ��05 �\�\�p��E�>@mځ.�!��	�s*JP��+J�zd�y 3쀀dʈ���;-��-9$(�b�Ψ*��C�hD�s�M�
��c%���y͜
~�.���oP�n��m�b�?��'&�L���GQ̨������H�*�-Qd�h�/7�X[�"O�9���b�P,ڲJӹ8�<RB��K�`*bՂm+�$��>�Gpb�z�Ά�#�=��D_;^�F��ȓHe1+��6PBh��"�d<�P� �B��`!�V1N`��I�\~�1+KC�I@�� 5������@��� ^PK�C�?�-�a��%�t�K�ZR���+O~ �E��N�P�;��)�!�Ę�J�ĉ0V��� �o��#��Y���'�!!��/rVyy�']J���	2R���@$o��'��΅)p�"� y�x {5�T%Hia~��0&�h��G"��A�WAǷ{����cj�/jU`@���?�t}�W`��y&���RF ��a�����'\hpA�iO).�Lh�r��L�d�
M�'TxPiN+*�\H���l�	-�=�@���aFkX���G��s˶�ɴ�:Y�fe��M�?dN:��'�\P`��%,�xv�� `�q�'�x�@�d�J�ځ �yb��K��yr��Y�`�sv� �<�K4G�+lD��Yu�ǔ0��
�'K�������V$n��D���y�VE�1䋹�y��
l�8أdD\ˮ������V,~�Į��}�FeÙwR؄�p��4�X)�d�I��3	�a���B&�N @��Q�F:kXƕ1DB�v��У�
�X}~���=O$�k��J(PЉ��Gx�L<�Aj;yi�j�*?�����\�'4XM#�/L�We��e���Db�=z�	a�
�@D�ȳ�K-���٧o�0v(�P	@H��|a{"��10X�� �O�bX� F R �yE^���dke
f2%@*�	���9���x����A�.fD
�Ƀ9K߀1A` $D�\�	�p$0��g��a���8��'d� 牺~^��Z ��w�n\ ��<��cY�("�`��w1�����D��u3C�i���'% �O��Ӓ 7x�T$���ʻ&�F|�a���GT�=ຝ)>�a�� ��t9��D�9qe̝�2��<ިy�U��= ���q����7ZVՂ�7k�:�O>�\B�"F�P}9��凌o��I���b���4z ��!
ƩW�n��DD�&��	��p�:E��yETD;��<��s��$M��ᙳ��-��[�"OF]c�/ù'B���Ě�  \y��k�7B��9%C��J��=��3=� M�����t��(�.Ί�pĆ��V0r�	�i��9��(mF.4��b�E!A�>	��l�5�v��$�_E6p���LO �[����|��d�t��J�b��a	�tC �CR�s�M�v����gOtZ��ȓ%�nTr���k��hل�[�-��Y�ȓ}�p���E� ��qF�Hj6Q�ȓ7����7d.D�T{@kE-p���ȓG�VD�S(�*��lC���(����W�:F$b���Y��̫��D��r�*yѷ)��:�L4��?9��D%�lY���=��dR�K}<9�}�Pe�'E��uH��� V"��C��S�<�K�x�j�(���)\rl���j�剄+@�P�1-��Sl��]X�%�.l��P�����V��Ɠf�6"�G�7�8tPA��Qux@�n#ft�ʓ&XV�y`�'o��	f���+޸���o:"0���ϓ/֨ɲPo�<f'��?dr���o���ܙB#H�Bȸ�
Oz� i�J��D3���3IZ�x�Ƒ|"��1MR�X�'���Ɏ���������H%nZVe����y�LZ���d�K_�^��9��W�JĴ�<G�Gg�g�ğ>�2�BU�[6�����!C5!��Oa]���S��x�H�@9J)�PV�l؟؀���3<�A0�e8U0�ڳG>D�X�2#�#�
�kV��y�1p��:D�X�P��m*vv+�?R"���	7D������H+�ψ0���WE*D��Sa�C�I@�R*D_�NM���(D�� $ĸ	�7`F|R�̳2�Qxw"O�:ů�:V��Xu&��q�"OD��A��+'^�9"�#
~.P1"O.��cM܄"eX@�t�Zw��(�"O���b#@(z͐�lD�!p���"O���ҫ�ƹY�h[-m@���"O��՝`G\�밧ܚBc�-b�"O
r��Ad
�à j2�"�"OVͫU,�Y2L�"¤=Ue�@��"O�%�́�Z����Y�T2J@�g"O��s�F- 0�\P@$�"Pd"w"OD�����'s��3���0���q"O��+���4Z�9saL(+���k�"O�b��<W�f���Mμ ��pJ�"ODiR�&n:��꣎F9��X�R"Ohq9�Oб[\,q��)w���W"Oxa@୓�C���pE�4*}(�"O���T�x��WlTS2=[""O�l	�h�OTx�*r��$���"O!���)���#;���g
�C�!�d�$#�����f��,?6<Æ���&�!��;I�V]i�e��,0xܺq�͇'�!�$�2sExq��e�tҨ��E˩y�!��ώR�����+Z%��Yk�O�v1!�d�I�`�R�z�v٧�ȅ7*!�DN�P�Xi3HR�Kc��( ┝;!��I��*!��:H��U�Ե&!�$�5D�b�;5��s�hl0ph�<U�!��<XM�a!e��}آ�)��<J�!�$��,�h��s���Wf��q"��2�!�d�a��� �xdP�g�'3�!�$�1Y��1h��P�2���[!򄝮$�B��ެs��� $ �!��ME�����4T��4�5C�"�!�dFw=�4XW���^?�y�L��!�d��:�B@�?N���5%�4E!��]7T&I���=���d�	xR!�D�#��,j�l�Vn�Y�1&LB!�DþxzXxjgHI�2S6q�$@Ɖw!�D��Q<Z�p����q6�8����!��3��ȢA�F�b&4qv,�t!�$�?n@R���F�Pa� ��)&�!��ɺ:+J$�g�M>NNB����\|!���=&�d���_��|��s�!�$�����2 ��^��m��k�!�@�Dv�L˔�X�gy����Z�v�!�D�&l �v�߫~y��Iw�\�@�!�dW�dy�- a��Q^X�3ӡƸd�!�<<A.������& �/	!�� �V����11���A/��!���s������yV���!�� dԜ���
�5i2�ɣ��\�!�}�`ݣ'K�&S�&-Ս�!��9Kॱ�i�4b8Fx���)!�S`\��
���4$/�2� _�#�!��-��FN�$7.�ڃ�4OC!�D�i��؂gH�V((�7i�8k�!��	�;�F�1� 9Z$��ʀ


`�!�$�ܢP��#�<8�{��N�b�!���hH^��$�,>������Qx!�A�?%��#�֍K��p�c
�vS!򤁚 )�l�%�i}���a�I#<R!򤖱9��L���qc�gd4!�䟘jS;6e֣m��h��`R�H�!�� ��X�
L�z�t!����|��cq"O��0lU5~ul�� g83�Qc�"O���TeC�=ePMٲh��2���"O�)aS�D	W��2�GW����t"O�3ɓY"��@��|��7"O��;D.ܫqPL���ζe~����"OJ�h�I׷ B�[u m���g"Oh�c�j����K �F� �0r"OV��4*�0'[�4��	�ZExp"O��;���7B�c-U�N0��"O|lj A<yJ��3��͉ob�"O�A��.8��#P%O��r""O��cwJM�/�RŢ�`�)u�2q�"O���N�[3��ao�7o����"O�Yく3��mJ���:1l,�"O�]���ل�*QW��"O��H#%0i��2P.
��8a��"OE1��LWx!hP� �:���"O���%)�63��aaFޛ%`R"OL-�J��d������	�a�"O)�0Gٝ(9p�	cZ�+�ACa"ON�Zu.��`��٩f�	:U���9�"O,u1��ޜ��8�ʯ��I2&"O`�3�ׄn-���q�ZMߚ��6"O~4s�ݩ3o\�ӆ�^��x��1"O�}H�B\�i"���E��T(.�r4"O�aӱDK<��L��IȊ���`"Ou!��ޤX �	
QH�*��Y"O�E�)3<i{���/$���a�"O	�h?� �	G��3 �rmQG"O~���ʆRft�[��0+�0I�"O�T�+'Kp�q�Ξ~S:�Ц"On1ؠBA'Q�b�x��E-iI�ta "O*�S��*NVƁ �ǅA8���?� �Iәh܈�I�)�3X��x�ȓ4�(� ����B�"eQ&�Z�iIP���d�,bd�+�� -�z�NX�ȓ{Қ�1�D;Et�����WzĄ�ʓl�l��%��zC"��&��C䉻2k:u����}���S��š˦C�I2yK�Ⱥ7G��]8����УV��C�0X$v<��JD�,bqӗ��h�C�	����[���)
����<D�hc��F�,g�q�ф+IH��s�'D���  �}��MS'G�@9�$d'D�d ��0���Wc�?���Dg:D��1��_�Y����
�k�:�!t 7D�Ps�LT%m6�@%��
$�hȃ��6D��R1!��,6�����G}$.�8�5D��1��J{X�`��Z����-D���H��8{^���_L��(�O��\&�X���	*�9�\5�ȓ�l�@wdT7Y���I�Fγ �D9�ȓ&�>��7,����Ae (/+t͆ȓk�`�
5dK<�f��Ō a���M�0�B���.@8`'iOb�\�ȓ	P�Bg�W(�9rp-;P����ȓ�Ԉi�o֬8u�	r�O�-@{,��2N��T�-V-�	�@�@��ȓ} ��gFBW�Mh�(
=GMP���Z>�D*%튱^֌�;�C�i�Ve�ȓr�8�#O�|`�c^5n����[�F}��Ù��Rq`L���B�xDi�gS�Xf6a�Wlحq{>��S�? z���,-�n��g��+R�f���"O�Ґ���x�X�G��(�L�E��3lO�QBa,�V�58S�8Fdt�U"O�u�C?G�ȗ�ѫWĈJ�"OK��@i��3�U� hN��y�+J0R���Ӂƽ$�H�8���1�y̈VK.�Y.\-�|l�‚�y��P�[��H�1���z��]�`D��y������ZejR(*g�\�bB��yrA�}CR9�LX�%�4IqwLD.�yBĕ�5�H�������g�<�y�O������	�h婖���y�A4A��lH��[?t}R��Ռ��ybL�-*D�n�h�zȻ�n��y���+1�>�iǇ 2��XƉ���y��Gl���	gP�U����Ά�y��4Ν2e*_�-yu*�y� �2Fg	ѡ �kΠM�T@���y��}� �,];��rd!�9�y�L�Uy���f):�f`p���y�
��(��(�M!��`j����y� �0��!+@ρQ�D)UJA��y�@�`N�T��#����
��7�yc�n�r���)�#L}�G��y�N��k�����D̩~��12���yr$�>7�������jI3��)�y2h�z�jy��D!̨	a��ybBL�*�N�`���&�l��$��y�NG>w�1q�A�#��`��o���y�"��:+s��#V�鲪S �y�ģ�ђՉհ"y�e�q����'D��٤�[�*ӎ@�^;���:�'�,�:�E�q[Xc��.+Tx��'�x�Ip�/3��U� lųLz���'P�Q���#/�l�s˕�LMD��'/L�Pc��3{�}�r�H�Wu:��'M��Ip��2`��*�]_$��	�'�t�F��W"j��J�5SѨ0[�'����i]�v"�0��w�D��'�Bw���}�pP3sc��{�'��tb���qU���II0hvƸ��'�Ba���@�&���'��ZʤH	���'"XYf�4k���!C�ص(Hݫ	�' ��Q7���t{vQ�B�2 �Ɣp	�'XN�X�/�#�(�BIh64��'�~�h����Om�,Hr���:��'�&��b�q�t�*BA8YZ4���'�.�y �4�Z�B�G��O�M�
�'��l%�$n_|S`S�0A���'�lh��ׇvN����)�4<��'fik�I�U#r̒�eC�}(@���c���He��TA�}��i�f6�Y�� �(M@��"���j�} 
��"O��c
�$
z��UjG�bL�{�"ONL� D(P_�)k�*H�y��@J"O��+�	 	�mHCɜ#)�hk&"O��5k�.,��ɰ�IU"X�C�"O0�Rth�$�f��?)
��C�"O
���	Q���J�Ϟ�I�i
d"O��xE�a��&ջXҚ��C��!?(!�d�Jt�ks��4fa�)T�/OC!�T#V)s4-Y @^�Ђ3��MU!�Br��0��V�f[������ "�!��W37�v��hE�4��	2��
/k!�� :,[�Í#cJ��wj�s�V��"ORm:�d�K�-�o*4�F�"O���3�1C�z�4� ^���"O���$'Y��IR��۲d`�a"O�+�]p��H�bˀ�Z�����"Op�{�$�$���q��� *�k4�yR��QJ�A@r�VLr	{3��*�ybj�$8#N�KX怕��K���y��]>��iR�MHVk�FG��y�"�-&�*"�8�i��	ŷ�y��W�n�lp��l�7���� i���yB�ֽA<��ӄ�*@=
��D�yM�Ud�1�(�&m��̟��y�,���\�U�D�D�x9bh��y��٨;R�l������!Hqj�'�y�7K��Zu�ԉͰ4	t�[;�y�¨bG�<Qs���~e��NB��yR.��$n�]���	Q2H��k�0�yb�T��*ܻ��>7.�:�(�y�G Z+A�!V+~H���M*�y��W+:�6-)�6�t�V.���yr@K��]
	�.H.���'��yb�S"B;1�lS���`��Y��y��ٺrL��ZG�F�4�ӂ�ӆ�y����>"���="S���p�R��y��/Y�fi��=���C$���y�	N���D��T����!��y���d�����fI7<�,L���̪�y�aWZ����f�6(R �@*I��yaO?��k�C���&m"! I;�y��F#z۲�G�N ~\��N�#�y��z�D³�Q�I}�%�A�Q��y��t��9����'P��l�0昡�y2�/#8�A�P�N�`mc�*�6�yr���34.'&�-t�:�00W��yb��/]S����n�~aaD���yb�t���W(i��%��	�y""Ϝ7�����	?I�Ԭk�Ꚇ�yB�:U�Xq��A�Uk�#�&�yR@�'k���F
 �6/~�*��I��y�AW�<͈���]����5���y��6Y$���f�!SP|��D��y�ߋ�n|q1%�N����!�y2Q2�ݡd�L�?�.1�V���yB�� P-i��ݴ/W��a*ڜ�y"�]�-~��R@ۀ-,�x
��J�yRB�	��W!�R#L(� (��ybjQ�k�(�K�	�6�2�pG�0�y"�0 L5�HZ4���jV�I(�y� �a�H�5 ʬ0�Y*��^?�y2��6'lu0��#�"tA��y" D,�ɐ�ٳ-�-A��>�y��ެb�j��� /�d�kF,X�yb�^�5�����5��A��y�i���4`�j������/�y�B�zhVU[5]/)�|#�B���yR�*_�HJ�6�� 1�n
�y�oӪb�rw��x>�X�JN�yb!��2�l�ʛ%jb��A�T��y�{uđ�b�ܸd�X ! �ó�y�G�#�P\ZT��
fm�� ��y�"���qĚ��9�W5�y�ě3@�6��Ԏ]z�X#T!��y�b܏Ulԥb�M�rvf��3O�(�y
� Pd2'B�>= d�q�͹:`t%+t"O�9�a@�-cȨԤѐ\A ��!"O��Q󩗊>��8	Uj�~�� �"O��"*V9HO�9�!�Z2?RzA%"O �(�0I��x��xFJ��'o6����ٯ��$1ub<�^��'�ιZ�솈s���r����p��r�'�R�;�&<Y@v�k�n;�'��͛�HT8,�Z��K�eE8���'uƜڑ-�s�p!X�FM1en��:�'-�4�j�tP^0"�d�`�L��'�!�Ê��� �K��  X��h�
�'m�(Rd�:��  χU� )I	�'����oŎ�8�SBCW�hT2	�'���Z7�=t<�C2�&��z	�'�������|����a�ֲ�R���'咭J񤞓F�+A�ߐ_R�l��'�ā�w�_'��ݪ���dJ���'yFZ����(�VE�0//>���'��Ī!ʀ%Q`���gW�!"X��'�	�S�Ҽ��)CT�ӹTxMJ�'T�	e��
�[��%D�zn�`�'Y���Ǆ��9\x��E.͟
��MH�'c�����Q(:&��eE@6E�'R��coڐ�BT�t�B5�J�!�'ol��ڵ���ٳ����c	�'�L 2v�H�~�>T#s�Y�$$����'I��h˜��TM��t�@�''P�R쎼�ƙ����wb�)�'�L١6�їgv�M��Y�f��'qhc��j�pr����J���K�'C"�!c*P�b�L9�ʜ/-�A��'ƕkEj�,o%X(Q�<5X�i�'H��y� ��C�,ăs��Z�� ��'�vZ�m 3��1(P�� d��'R�Ѓ�%�#�j���� P�1�	�'*�T�î���R�C������'$�`��L;=�N�8w�GK2��B�'�̵��bg+��q1�'Dq��y
�'�tArmC��XsP����Q"�'3�Q�F�� 5��J�C�ך,�	�'`�l��	�.���L�&w�
�'V�Q���-��ٺGNf��!��'e���ë����eQ)�h��'����i�*Q�� צ��6f�I�'߼�bF�ΓcA�E�S�?_k��z�'����=B1��4$
[8H��'֤Hw��U�P\��ƪ=���k�'l<�s�>2s����*ԧ5j��'Wx ���[:3b&����'+�(��'�~Q��d�7LFJ��@���!)��'=d4�ߊn�dPOݯ}���':ܔ�2`�#0�IW �
x-�	2�'B�1J!KE�T�F�XcCH#�����'C~���� ��mcJB�{nh��
�'���Y�"��DQH�?(Zh
�'�ñ�B�)(�J�Fӥ0���	�' x�z�O�R-B�U -ha��'� k����=k���!�<KKJ��'���K��˝$�D��ef��B�`��
�'K|�������`�e�ҋ:
�B
�'؍i�CB2(6,<r��6N�R	�'X�Yi5.
`�I�a�1�6��'E�d�:yq�C�K6-f��b��� J��v�"T�^e�s�Jc���1B"O0�����q1�����ؓK�N�x�"O&�P�D�_����F�v���id"OR��0��?.�H\��.��xg���B"O�����n]j
7��u\�pi�"O,��5!��Qh�+Q�P�H��"O:,s��0P�ܸ����@2-R�"O.E;V�q��<��Ë=T��"O���j�9�@�#���M����"Oxݚ���D���8s�^ [0<�+�"O&�괄V��J�8ad���$E�"O0}j�L�F��k�/���S�"O``��d�8`8�֡�9=��8 "O�y;����$�� ��#���jC"OB-9�'c��d��D���""ObL*�J�[���d���<)["O&�Ta٨,�b$� ��x��Y�"O�;���M���)��\���=��"O�7��E�ndRO
$P�"Q�"O�����L�g��A p�F�`���"O�8�%�6"�"�&NX̘IT"OB��'E�U>�A�V�r>�mx�"OX0i�˖'d��1��cX�R/B P�"O���g�8D۪)��ͥA(\��"O�Dx%��6��)�r����\"O��[��Ш �� ��%��� �5"O-s��NU������%b�{�"OB%�#n��>1�9�c���h���#E"O>��l	�b,��(��Yʶ��"O"d�JJ�}�"M{�k�x�:�"O�H��Ùje u�â�&6���8�"O���i�"rez��P�J�1w�́ "O��1���|U�V��
�k�"Ol��	�n����%�:F4 �d"OH���X�� H�s擋( $H�"Ot{�aH�id��`��5q���C"O�d���6;�l��I��.d8��""O��s"*̀$_�T�dV�y'n���"O��B��KSN�) ��9sp���"O��Z��#|궘��-)S�,qe"OAQu�ê3+� `�Z�3M6�("O.��6�P�8����^�k��;�"O2�cB��J�<��eJ}d��F"Ox���N)ޔ�҃�C�s���"O(�+�˛'Ԙ���X/o��5"O���G�%�:d2��2R ܌��"OX���ӻ1��H�E��5/lb$"O���@_�s�����"�0O�|���"O~,طm�uT�(��X�0N�q��"OY��`�d��b� f�(r"O����IȒ/���j���jx"Ob8CpJ���yY �65͚���"OPX�E�<%f b�ϋ�D�N!Z7"O΅��n*�
S�Ǡ|�|:a"O�݁b���Vj5��޶���9�"O����Q�1�,(g+S"��\��"OX@�f&Q���8���}2y�0"Oh���&PlSB�$�0Oc
y�7"O�HvE޾g���q�=d���P�"O��QDZ��p1�!��D�l� �"O$mP �,<�E��i�P�,���"O���f��8Ǫ���>�F4bw��j>M+o�az�1�U�^}R-K�6D�!OE\kt�Cv @/z$|A2 �5D�� �L���]`J���ߵ�z�+D"O���&.E7t��(r�ʈ�i�v��"Oу�@�f��f�K�a>��k�"O�I�Q y�� ��"��6;8�2E"O���d鎳b.���^vZ�QW"O���̕��b]+B؈��"O���U_DӐʀ�(M^ �%"O�xكL��Xub�Z�)��ge����"O��c5��#R�6��Ĥ(�f��f"OH��� �n�d�d�
�D�t��c"OT�w� �z}r=���M�.��"O��@c
@3�s�X��L���"O��P�-{iN�"�ҡ�D<ɒ"O���ɔ�(5��HX�K����a"OT`����	R�M�aD��n�)s"O~��fJ��J�&�[0�:�����"Ol�*��Ȗa����q׶o�����"O��c(�)�C>�B�"OZl)b�Fd����-��$�s�"On����F�@�X3��УP���"O��)�g�K�d���G�ԛ�y2#�7)�p��-�g��i2@9�yN�_��8�3�0D �P�M��y��H����m>2`���'�޹�y�!C0n%�(���ɠ$�0�@W�R�yҊ4����`���s���k�� �yRF9բ���֏n˜��퓃�y"fÛa;���$@�<T�dJ�D\��y�G˻W�x]cB&S8��*r�ߎ�y2���0����	B�2JB��R
��y"-ж@��Q�d��!.a�M!e�3�yDYG<q�b6w�������y2υk�X�Ci>��]"�����y�'Ի�n#w/29O��{��;�ybj����*b��:.���
�(D-�y£�*�X��w�֓.��P��$�"�y�ɛ8"��y�@N�#��!�T(�y�FE������3��m�]��yB�T��}���9$��j��ğ�y",�-8ʉ�䖓*�>):f�F��y2�_8;�RyuG�k�����ڞ��=�O��`pT�lhv8�U�QY
4X�"O��a�Q�<cDx�4�� 7l��"O�l���đ
�����1*1��"OL�6�_�,R0�P�ѵ'�9�"O1"���U\�hf&��Z��"T"Oj<B5�N\L��ەM�v�����"O��R#�dezqr�NބI�@D��"O�!@KƎ4`N��C�рd�rH�"O��0��Ɣ7��傄!�V���)r"O����j_6t�4Ps�@�0)d��"O.3��T_�1�P��OM��33"O�XF��Dw&4�͕�FӔ��"O��ȥ�Z�YSD��,	x�q�"Ob4K q%h��
3#�`�a�H�<iu�R8��Y��קB�#�B@]�<!V�V� ���V��$w�pi�Ώm�<�sK�.@�@�A��"ZB̍�1�~�<9��}C�}i��@�DeN���I{�<@匢;�3`�C���4�Om�<)��' ����2ʑ�0Ș���BN�<Y��@���j���Bh��N�<�3L�iB�QХ	��RI Pq�`�<�/ެ^[�`���Ʊ=��$a�.�^�<� M8�����JЁ�ꈱZ
�x��"O&��r�W���k�ɍ#O�8�1B"O�eX�ÝIPH �q��'C����"�|��))�������V������':B�	6���K2��?j| �)�E۴n�xB�� +X�p��ݔ:�� AM��<NB�ɭvl���'B��DX֯U
qnFB�Ik	^y�1݆gMn���NG�3B��8<�"�9��z���4��A��B��>
�R`е @�NFT�J��fC��&Rb�u�RJ�"& s�
ܸs0��?���� y(�j��Q0`k�%�D�y�!��oen0�����j�ڭ�� �{�!���oV��T�P%(U��C�!b�!�D25���p`��Qh�����3��'�ў�>��W)=w��qʟ�D5<��A�4D�P("[/:������5\Y�7�7��*�Sܧ(M��c��n�`p$&\Ȃ0��
U�������=�ɐ�1i��j���r�MZ0��s�m�6���ȓV�N �A�W�Z%�dK�o֮[Ř%�ȓJA���#*H0�23��D �L���T!.L)��R�(Q�e�O;����ȓ0�F���-(<j��K�:g��ȓm!��eY2��@��T�/�̆ȓ:��
Ҁ��N�$Q#�P$R%���ȓh���CǏTM �������Y�� �PL���A���3&	=rj��ȓ:E�وg�ŊJn�u�G	��LTP|�ȓ�Ԙ9c�m������7��dpA���ҒRx�ђ��Vh���\ߎ�ۣÁ���]f"��	�B��!$au �x�*�Y��q�ȓ-	`�����>Q{|)(�cR81L����+�ܤ�r�(5��B�ӵ6�V���P�pPzР��&Ҟ�#�1�zp�ȓ ��8�����h�HB^	�~��ȓU�N��Cc�"`�`l%�W:���ȓ6<vm:ec��PX�Q�Y�ȓ(�u�4jҲU��t�&X�ȓe�V�Kr��f�=�c��>-��ȓ69Z�u��=<��P�2N�a�Z��ȓf�uz�dRO�09qD�Ve����ȓ�JPH�b���n`I�.O9 ��ȓ4�Ԁ��h�1�r��D��Q����d:&y���=m�f�4��8*��m�ȓ#�V��BD��4 |�-Y�H����=��7哌�>�E�^9/^8��Z��9CF�#Vt�8�J�	�ć�2�>4�Q��!<�%Xf�7i\Jd��S�6�!TMT(}n��`�w�f|��^>�쓵FA�
[���g��� ��q�ڼ"�a]
1n�r�EԊ?���ȓ��p�h���R�)��L�\�e��N���SG���{a#3GX���"%D�qqW�v�`;���/8@f��#b��H
=4+X$����k��%���	JyR�0[)�	�W�l�#�AVժB�I�[�2�
�㗔5lB�ir��.ՒB�:b<���Z2F�,�X  �	#J"B�I��T���we���b
O�;�C�	G�Aj� ��X�\#g�ٯ#/�C�	�r��[�b�>HL�� '�?=�C䉵V�,��J�j��p0�e�*g^�O��D�O4���� ��ZG ��^:%�1g�*��,Kf"OTl)��*T�T�X�v�6W����6g>t1��P8Q����QN-�B䉍1�H ���׳լuH%�f��C�	�;Fdpȧ�ԳSI��s@���\�C�I�d���2�Z�"$#�,�7:��B�ɷ2���f�� ��M؆�
�	���?aN>���I� ((ex�K�l�� Ă7?!�d��=�b���1���CA�%<!�Y'X[��ʳ���*���!���<Y��P*�2�niI��P�!�!�^-J˞ 0H� $�����#�1t!��9֞ЩďU7�$=�e�ל4k!��I&�yip��kn>�!�Y
��Iv�Ո�h���K�^<j�R1'!|p\0�"O�mS�"�""�6h7Kq��{�"OP�A��!?�H�����]T\��"O^i�#A�����ݦW�V"ON@hf�����K�DF�[1
-a"O����'Y"�i:Vn�!"���C"O!��#u��VK�P�r��|��'�0��!j�/4y
��|[��8���xr�G�o�rXQ�Ѭ,ǲ�vG�-�ybN B�!�i"(4&���4�y��8���ZP��V����g�*�y�ԫ!�j��eM�Mb�}�W�D��yR��5�F@p��H}����LB$�y�lNi��5���rcH%�f����hO���隥!]8(����!����\$!��n��%���/"̈L����|!�䞐?��0Èn�,�x���;9!�Ѭf��a��Ŗ�h�@�� ��J!��/N
����*��Qh�] !�d��P4� C�����ęI�!�$�/bJF=`fꊡp���Z�V�!�Y�%��0ڗ#Х6��cd�դ4c!�ݠ(o�5a7�TC}BlD�K�Vx!�d�lRX �I�/.��|����'n!�$C�vMX�pG(��)��D�Q�D�o�!�ίI��Ɇ��{�l���⛮)!��[V���@�M&X��"��(�!��7d: �p�Q�v?`�a&�
z�ўX��Sm�)2�i�X�\����ѤtJC�I�g��;��̍(Gx��p�9A��B�I�j����0:�X�*ãe������d��fC�;��p��O��h���{�&�a���Z�T����eW"��ȓԌ�%ԩ�$�#��X6;h�m�ȓh������tbuc 5���?����0|r��@/w�x��H� h��ivF�X�<��� ������lFyY�D�m�<yք�$F��*���[����G�R�<�"d�/B5 ��A��e�P`�J�<��֞�葲#cN������]C�<��F�"D�EZᙼ!?�Ǫ�@�<�@@��=P��Ӯ��"��e�<A� =2P@'N�!���c�l�<�P�ſ]�.1cl��ă��3D�4+�懑zRYk���39pqi��$D����-�+U�	�i�P^]��H D���%�-
lhj���sf�#n=D���W"��v�n5���7M�T���@:D�L1�Ƈ���d�!���&��.D� Cr��5^t5�f�8x�>�Rn,D�� �X�ME�j������\#�TB�"O�t2��H�Q�TR���48�� WX�����>5���#s �<��xJd�_$(��C�	t���c�<5�@R���,�\B䉒K�v��h�7�)c�\�[DL��-?	� W�&�^ R'�Y�v�*QK�oE���̓jd��m r�r��I;&$Q��p�~��QA�<;i"�.�4;�V������� *�u�Pp�BU.�j�ȓ B�t��&��
x=0iU�p���ȓo8�=��gb�E�I�����]����ȓ��Z� '.N#�X�Ɠ\I* ���1��I�kԈQ�������hO�'Rΐda��I�O�������Q.q'�(F{�����HB��F�;88z�&F�y��A�@�M�P,Ƃ�!��=�y��:��
�lʢ(cbƷ�yrf�.Z��vH�^5��(���y2�R�NL��B0H>j ])p����?��f&�֌٭S�,0��:rA��*O����>\2r=Y�*o��W쉂�!��D%�F�P� -�qj�4:�!�$;R�d���].抹��. !�D�~��q���U�N9N0�`�X�!�D�&1|<)h!bz�$�{6��%NL!���0|���Ӆ�0E�dY��w=���'�L<H��ʖ-���3�a�<�T`:F�'�!��@!T4��i�n�,9�LӯN��yr�	)�������:s��e-ҔAڒO���D^�*�HH��@� ��� �\�]b!�D��:��DX�*�Fu^!�G�$�!�d>*!sm�Njb�!c�Z!Q�!�Ď�L��*A�ެQ^�8c�n�7g}!�D�l-��K�iL5�i�n��u�!�jC�ܻ�Oo��z7�
+T��}����`��Ѳ\��&<ƼQ;��O~�=E�48D0�b6�ɾq����B�4�!򄙅(	��&�
Y4�1�,Q8 �!�$ЛFDa�" s���� �-@`!�����>��x8UA�D��č�|�v{�
Q�DnM���A-Ez`��:�	�D�p�B���n���J���'2 ZC�I�$l�*��>���C��ߘ]�C�21�p���[�ȹ��_�n�C�I+5�8<�A�p^ R���4W�B�Ƀ`�X]`uc/r��J-M�B䉋q2*hcU���@�5C�t*�B�IV�1�ḛ&�| ��S�T�ȓ*K�,
��~�>�RՊ�PԂ��z-���b ��jZ�.L=\)���?�ӓXe�1�QI�:n�*9ʅ+۵@�L�ȓ[�h�!Ʋ7���hU�ԥ��=�����kS��z�iR^,�ȓK������]8\�
��2�L=��I����<�� �5t�J|1�$bk|a��EM�<!q/J5o��{��6S>�E��os�<A!F�.Hq��c�	O�MQdKx�<���X����隌�L� �M�<օ�k]��UC�M�:�#��~�<I�f�.!����mҽ6
��cb�x�<�@a̗M�4�Ë7i/��Jj��<ir��#{v M+��7m
2�2'�|�<��˔'���i�'�2x�V���L����e-�xP����G�f=��&A$tnb��S�? \�p�~�xM��p���"O,�u��T�UAA��O/z�H�"O`����x`�8����/KlŁ"O��A���T �R0oa�"Oz�Ʌ!��BEU:ݺ��R%ف(|!��ߏC.�����q�M;���%R!�dܝM%��a$#�li�gm�yr�'���'��V>���r�ƨ��bU�5��ݢwL�!F��ȓi��
`C�V�"`�Hψ
��l��$,"���͝(ݦ�s�	ه-��`��ws4��AIkh2�P!�/It�i��#z�����~h\�+.~`B�I�6
�������U���G�NB�ɟ� ��Saǆ��y�E*�	�$�Oh�$�O���|r��'S��r�Ռ:�e27��$(�رs�'jPm� �x�d��&aB�'vJ��B�'�ax��q-vP:�@ٸc���[�.��y򫔮e�z��v��?`�0w!�yr%C��C����X<���9�y��:3��-Ŕ"����C��yr%�v�0M(oĸXt�FV�?i��?���?���?����vs�Y�TO�ZVKe��%�1i�'2�ݹƣW�9��anߎj�K>��,&���+L�7l�Cs��H��a��-2����/,��r��%}f��	 �]�v�X��JI�o?l����	K����.���a
7�Mk&��:
��P*O��Hp�Y�!W!RU�H�z���A"Ov��F��\�\M��f-q�a�""O�,���Ƚd�`Q#�ğ/R�88����F�t�Kʳ����H:B�ثL4D�<@��S>`��jɌp��pF8|O4b��
 ƨ7GN�v�H�en��@��<���S��2�9�Ӿ~ $����z�VC䉓	HD�� `��V�ָ2��;.��&@� ��J��a�/��M ��ȓhp �b�'��}�0ppd/�2&p9��|y�|ʟqO�$� ��d��MB@n��=����ȓ3YX�Yt��3ƕ��VO���al�p4lߠ]�,(ᑁJ�r4D�'�2��<�A�f�S�8�m�sa�(~��C�I9[��5���B�F�L�1�`I+V� �O�O��1��9f�F�Z.J��鳦b�)�HU��m �1{a5U�t���Mܐ2��	�If�����upŠ`,0��Ð�24n�ra+(D�`dF1/B�ak��Q*{� ȓ!#D� ��C��2���-�b��O���2�)�'�c3��-X}�X�GI�8sF�(
�'P�}
�N�B'����m��6>��j����O<"|�0�KU�(h�&Ç�QXJAq%�M�<�'Ljȣ6ꊋ$��d�GyR�'�OQ>��!$I�AȑX!G]��u���!D��Z�G��S&��5�^26��a�'�=�O��]v�����m?�t�&$A�g{�����?a����ׂG��y�afU��	1��-��C�I��M�@��6jd1��թzТC�	8=�,�"	�$�lp#�x���G{J?}	������Br,�I8~�Z��8��"�Sܧn,����EF�<����H���ȓI��tQ������x8� /�84�ȓ=wpl/y]tT(�h��W�"p�Т5ړ�0<q5��+�iEE��0��;P�p�<��� S���
D)I�8�\����a�<I��/̀���uΘU{��S`�<� ၱ���1��Z�R?W@�i��|��)�Sv����R�>��6@L�l>�B�I�n�d[�	J>x��!��5�vB����)3t�O�f {(�R�C䉪0Ո`zV`d�>|�T�V��B�	�\��CE΋
:���P@�ڝ��B�I�<!����o�b������1�B�I�"�����gR.hD����T�&ĒOH�=�}
�&\|��q@��5JB1�ϋI�<�«߂cT&Q�Ǆ(K`F�Yd,�H�<�2g̏4Xܔ��X<��9�R��D�<��^�:n�h`gKǑp���$��[�<���1Gfi+L�	�\�� 
FV�<q�G�a��=C�/ �T���Q�<�uE�$�bd����_��]df�F�Ij���OU2}��2P��@Җ�.�!��'�f����*p����cL+;���'�N���-��|Y����Y��4��'� ��DN̸��$:�֞KF�хʓ{�h��*��F%Rq#����ȓ-���1*��V�D(2�M�)�%�ȓm�0`P��6*���\4W�쀅ȓs��bď��ru|"6/ר"�h݆�<�1A��3M���%O�v��!�ʓN�c����F��<�� ��B�ɕU�ʕ�'/�-.���#�oM;��B�IC;XY)S��`� �;���#?�E�'!��'������R�0�wŞ�(���9	�'eP| ��L,J��9Fz���"D�p"W�\27��8�ǖ�>PT��%;D��тD�.B�nI"��l[H\(�/:D����[��(�hK&x�g-D�adJ��4jZ>-Xu��/9�������I;& pHT���A�:�ۗ��up�ʓ�?I��c�޽,��-�D�Ս}�*��ȓ����Nݹ2���92��-��\��p���C1fڈj�h�Q��ʳ�(؆�kI���4KڎM7��[h26M����,~�!
���N�LlC孟,�v���<Ԭ����$8��yw- H�@�'��'Aaxr/��.�A� !a��9Y�E���yK��(�-��^rL{�Aׁ�yBD8q.`��)�Gb q`�I�y2��|$.٥�=�^��G��8�yR�	/GMP�A�)J7!��+�C��yb���3"�P3��(p(I�Ɩ�yB={�9��\��@h�Z�䓋?ӓC
�1� �X�=����V=��x��죱.��]���+$N|����F��!؃��+B��e�;8��ȓp�F9���^;.]a��w�lЄ�v�j��B�*��E2Oz��ȓ3���FB�:-x� ���13Jp!��(�\0��(@�0Q�
�	݇ȓw\� ���7��1(bҜ(h4Y��=^`h3S�KfN��LGt�*݆�ZZ�0kF��H�/.OV%��q���D@��:��r��,2SF��ȓD��hVnA(u}�] ���-Thܡ��Y�	2�M�Q�|}�ԩ�0MBx���96ty�b3�!��h�*6U��cy�H��	��l+�����2d���!5�����U�o��`@ӌO�乆ȓe��Y�l B�T<�F�=v�І�S�? Lī�ƿa=̬[�.�w T�B"O��bA��KN�9s`�[�x�W"O �U%P�N�ֈBEI�;=HV���|��)�0s���Ua) �d*E?&�B��7V�����J	H�ĈXF |3HB�I�rߊe��H@�n����e˶c8~C��+1�5���:i2bjwE��v�vC�	$ ���CՊ\\F� H�)mwB�I��6�RF�efZ������`�4C�ID�8`)Ƅ �h���m�C�ɜI��ReċZ� hCdݴR�C�6zfȩ�thO�p �����2 �0B䉟qːI��բ!��ź�ǃ��C�2ig�)�&$M�KV��
G��C��
�	+HX�J�ك,c)�'?D�Bgh-��P���U�a��ʔ�=D�D�u`�K��[���6(:����D:D���g��U� Հ��N�Z~�T7D�bs,�4?�y�@fW�b1Bq0���<Y����(�&�I�u%<�($h��C<�1�"O>��3��5\�Ԫ�H��"n}�r"O|�P��$U��QQ�&Ѵ�&Ms�"Oxa���n8DE���;.�����"O��Xd�� T��I��?���c�"O�B6�J8����͌V����"O*!`�J=0���Iţ��~�Y��';�럼����Y�r�Q?�f�Sc�
hۖEz&�,D�؉ 
ۮ.r8c��ZT�Z@H7D���矗�0H+��(#Kp�+��)D��ˢ)�/	T>��Z�l�Ph[�}B!���k�01�UxS���E�>2!��?v�^HP`�4���6@�
!�%.�4��A,,���F3l-�}��'�$�G�`!���.����0z&!�DD�w��x��M�w�`SB��!�$����+pn��_�r����~}!�d��x�茱sc�Kwh9s�B��!�$ T}��ȓ8��٣���R�!����S�F�I��p��5f�!�dֵQ/�U
`�0}�}���Dvў��?����yS=o6����999��0�A+�?��'U� ;�BW4Zx^�I�J�~3L���'��0֢Z�79�!0b� 	}W>���'�NP�m���A��U:i���y�&y(BI�"6[)D�3��֔�y��̛,y ���'F�p����yr�9gi�����;6���	�����?���t��aO
�ia�g��tt�Y`-O�����h\��eK׉I��CD(3!�$��P�D��7:��}3t����!���\,��؇Q� Mٖ��?Ha!�d�c��Q��WK�YkUN��N9!�$�R�}�TnX9�L�R2-:*!�]"�����&=���+s
̓|!򄜯+��)��J, �"!q���� |!��8&:���E�@�׺�yiÝ(r!�d!:�a�t�� �8 �g���!��1tRI�1����[pX Ɂ"O�*��߹nL���`W6R���B5"Oz}{'�� 2����*S�C���#"O��Q%�Ir���"5�_�V����Q"O��[�@��~{���E��x�<:�"OF`4��zvA��F�LfF�C�"Ođ#�ݡ0�p��J�Y�5s�"O� ��$�s�̅���M�B�:�z1"O�Ⱥ�H
e�N!7��Kc"O4%ZQ���Һ�v�?	lڍ�"O0�8����S��)��=\� ��S�|��'��e�t�	}0\� "̞Ȕ�'ABU�ׅԝ22�E����
~Tj�'�B�9��i��,�e

K�l5��'5���@P�
�P��͚H.��'+���D!_�_�l1�bԳK1�59�'.�8j����]M�R��H2=���'FH|�sb�/U�J�R�C�����?9��D�O�b�����
bx�-(�́�^�ƔA�l�O�C�I,2-�N����Y�U���
 C�I	@^td
�*�.�1�B�
#��C䉃K�v@8��DJt,���AP`C�I�6��șQʘ�<����l>C�I���%G�C�堂I�,�
C�	xh�ǋ=^Z��A@^�`�����O�=�����)���'��e�Ek�(��}p+Oj�d8�Od9i7�G\�A򉘬)	�Ih�'��\�����h��4R��0s9����'���#����^�<�g7xx
�'��d�A��v�H�VA֯fZ�8�'o�!�-(���\�[8�H�$�#"���7�Ȍk�\��Qʜ!�!�DȘEb~���"�*���a'B�Y��'�a|��1\<�SRm�6_�ĩ�5����y��cu�ř�l�h%nх�y�d�#0�ްClŒ{�%x˔�y(̔��%�ej��j@F��0�W!�yb+�I�H0�%*`�J�����=9����$لP����Y�EF�E�n�t�!�P%gT\��u J��'��&�!�$�25`��0D�'bEK�ԧnx!�D�2O���#g���_@�*�D#4:!�@�?�¨1��Êqd�z�ƻ4!�ě�,�X%Án�@�r3A2J�!�D��M���8�I��6��Yʰ@�+1��}"�'�b�'�P�KsiA�o�ā����pm!�d�s������� V�����5I!���OY�T�C.�#S��Q�ŕr�!򤄹w�����;~�<hz��6:�!��$?`��q}�h�"䌰~�!�T�b�>�����EL
�z4�׉U[!�$E*n��'�	V�X�zP�ߓu`��>Ol��%��R��v���$k�z��)<O�HS�$��sJi��A�v;X���)D��t��y��S7���>�@�=D�<d��9[�Dib��0Z�	�`6D�p�g�Ԟ#��c�U
���5D�D�W�ι*������	?>�[To5D��9���)���BR͑;3���RR�/��0|�&m�.��9�-KO�zU�K^h<��) /YDMIoL$6,;vN���y��Wӈ��A�%24�P��&�y�a�?����c@�����
�
�y�I?T�e��� ������y�!�a��aG�:��r�!��o>����3��Ą�{'�'O�=Of,�a�))��p�0N(2�H<y��X>�˂m�k3�lH�k��P��G�O���0>)P"��i�MY&�v]n�����Z�<�#�۱dsJ�!�#�5V����s(S�<���F�\>��ֳM�;%%NN�<� �H�GO|nf�8���?	�x��F"O 	P�ŉ���H � o]���'ў�I�'ovA�!��
P��5��[Z���'Zd%��gB
f�����
Pn�3/O$���6^��� %F��u;
�'�~s!�Ͳ9���K�7I@	3e�S!�Dμ;��5�Qd@� �(��6��"�!�$�.*�8{6L^7~"h�ʒ��(y!��C38�4�4���cr�#��|d�{�\�@ur1��>f�Q[��L<!򄍨cښu�d��9Q[����"U�!�$�?�z�+F�[>��R��·(:!�ą!ddEX5jO$���S�ƒ�!�dХ`B���C͓w~(%ѐ���5!�3���Ç�{�iHE�ϒ@�!�$1@�<��I
<^
J� I�G��{��'�I�e*p��R�$x�!r2�Ќ[h�C��laB��y�����ĝA�C䉓 ���c�np�Y����-�B�		v���rjč`?x���):��C��R��t����]�^P&�&'�C�I�/���X�H%�"^�za8B�I;�iH����w5Xo[�*	.B�Ƀs�N����S�iZ���(e .C�I/w���d���T�$[���4��C�	4-��@���fY�z��+NܸC�Id�6% ��زA��T3��S-+.�C�I�7҈r"��>��A��;qjnC�IY��Y��o�%_�Lm�%H�=Oc�B䉄o�d@d�Z�N�^�aS.1HC�)'|���;t�x���7|�\C�28K��Ң�[#�v5!���v�B�	�󮁙�V#$Z�)�OΗs�*B�ɦ w���J��`sn5�$�A&�B�;I4}�2aU������+E�B�	�x�nU��&�M���rB��t�B䉥6����n��A�Ȭ��,�ckHB�)a�ȪÅ�XiT;b�� LZ$B�-`�x�m�we~�ӂ�E*C�I�	KD}:��ٽ-B�ѓ#L�B�ɿUm�]�� �M�l���t,�B䉚uy�!�C͍�a�c���]��B�Ɇ6W��h �ؿX���xEIҹ�bB䉘�P��H�"E������$VRB�	���iRƗ
%]��aGه-G0B�	�F5��%!Ԙ*�TH
��҈0�C�
4)rl[�F�0�rؐ�'N2��C�0h\)�č	0~��\ �9x6�C��e��t:V�оP��L������'.D��;��I!L.x���(��'ƈ�`�k*D� ��B[8<�.
Y2H�XjX��yÙK����BM��0 Q5Ϧ�yr�B�d)V��A�®?���Q�����y��?g��Y`S��#@@}Ac�å�y"&^(��\�a Ģ;�i�� �yR��2^�j}����>"z�$���y��@�L��0hפ ����Q��y�
O	3%ĸ�B�^�\�Ac���y҂PX��ɜ8^䕰Jդ�y2c�)]<�Hq��TQ���5�yB�ίO��!�I$&�	� F%�yRc
������!fP���(�y"�;R�x�uI޷\)h�A'��y"�ɛ����`˒X�z�!�aܘ�y
� }	�Bz��X��,2p ""OZA��(��Div�Țw���k�"O`}��-��SA��XS�}��"O���Ԏ@3~�T�G�;���q"O|m÷l%t���xM߆rSr��B"O�U��CM
%-����AӉ8Md�b�"O@H&�X>~ <(p��E&��"O\�FMB�Y*H\J�!^9��"O�]
���X�B/�gt�д"O����jچB��-��c+! �a�"O���鏊R��s�,ΗB��(e"O��;$cK/pF&��C�rު��S"O��i�����	0"k�8[�RI3�"O\yB%� j�ѐ"�y��K3(:D�D�  6X�ι�A��J�q��7D��0c�Xw��	��eZ&D�x�� D�8s/N�����I�7\^\iE�*D���R��3/g~x `��9>c�&&D���p0���5HڼU���%D����f�0�=�e� %3�1
��#D�0���.SC��Ak�%A��4D����^1
�НCD���wc|��#�2D�d��IK�b>�����c| �C�`2D��f& �"aG��:�e��0D� �h�8&��A2bBN"^H��p4-D���2G9��r�"΀8�Ҝ�`�%D��uh?{T�ɑT��!��UÁ�"D��B�^L����%L�# ���<D�6�W/%O�$��L�BKĘ�#Y{�<9���25�̚d�@�:ь�fOu�<��i��D�R��*?���P��I�<�������k_,X��,�v(�]�<)��˷�"1��A[�dg��(T�B[�<)�#��R�Fqk�������0�NZ�<��F̀CG����= A���,K�<�`a\aHxx�`_9bX����{�<a�ᒊQEp81��¶E^�!�I}�<Q�����S�
/4���@y�<i�N6Z=�!s�%3<:��Zd�_K�<�ǣA�~Ȕ#DM�(:U a��gVJ�<�#��s�Gߦ2�@|a �Fb�<o���ACP������A��Z�<9�L��Q�d���J�|�E��Y�<1C�m�R�,�\�A���L�2�ȓu���Z��Ԁ�J��O��jɒل�傽�e`A9}�H����|\ ��ȓ\�4ecP�I;3���P%��;!	��><� �'�R�6k�(��&�i� q�ȓl���P���<���I�'֋	b*��2�nq"�@�.jR�����llI��j�R�z����'�i��[3��Մ�S�JH�b�^#9�|D�"�Oy.�ȓN���ХW��\�`N�=���ȓ3�Z�h�M�"g�2U9t��7�2h�ȓKL�)kK��W��!q���}��|�ȓ&�$�	6�jx`�.
�<XF���#S^ (4��ps���EJRR�Յȓ~�����G�^m�&	K�����61���S��"苐�A�*����`����n�	���`E;]���ȓA�^��DR�J�R}â�O�;���{�>!1�cR7,�(M;�Ή��>�ȓ3�������-æd1�B�:�&��ȓT��}�F�� �R��%|��|��S�? "��([#3V���U'@�"O^|��%�EЖ� 1�T�\I+�"Od `��	�~�ڠx�ĝB�`A�"OrR7жV^���Cn�JB����"O>�i���B����glQ:<��j�"OPqgq�<A��*G$�J�"O>�J7&_�+z�Q(�*�6؀v"Or��aMG?����Q�[ꕫ�"Od�M�I�P`럒%���;�"O.)8aHLH��
k7F:`0�"O�%x�̬{TTyY��ƟJ:̙��"O�a�@�Q6���t� "%[`"O�+� W�=B�pJ�G���@�Q"O�L"�F�4����f6y�ܙ��"O`���+^.G����f�6���"OЅa!e
^��8�%��*�Y t"O�xQ!�W� ⦉�G$jd1�"O�l���(SJ��qB�&:��0"O�q�֥�T���k��	�|��"O�%��I���x 3��7��x��"O�y2S�G��yC�_$���"O�4K�����a�1R�ִ�B"Of�fd!<dx��)�R��q"O<�`� S� ~$�!�'G!6�$@�"O��X#(�0s�}����,��A�S"O��"��	jW	X!C�N���$"O�豆�,��Ӂ��h��f"O0�7��M�8ڲ�����<�F"O��r�*� �c�F�.a�H#"OĜ9�BW0t�9��� 5Up�8�"O��3&J��^bHI�ЌoXD�c"O�����ƒr��,WD݄Y�"Of�����M�l���DW
xh���"O�0J�+!^�%1C�:B�!�$�#vX�Z`��12���E��#�!�9M�ҩ���׈K�$4
�$�!�$��d<$+ c҄L��$C��[�4�!�ٮ ���c�مn�T	��A�\�!�d�qaXx�� V��iF����!򄜳lT����'@4p:b͡�\��!�$6f�bd�S��V#N-kpΎn�!���L��n��#�v���!��	�C�BـB�;0����y�<10��Qd��A��^º�&H�r�<ч�^!g� �;�+V�xބ)1f�H�<) %���1⦚�A���X�#F�<����%Q찰x�{<v-9�B�I��$y����%PL4����&^��C�	7�P�c$�YWĥ ��	I�
B�	�a&٘��WI�ځ�.,R<C䉡|���+��'�\��   R���hO�>eölI�qa��)���Ȇp�׮:D���鍪�������A�P԰�5D��GoJ�m����&�O<|J^��V�/D�8��#
�qI0]`�B͒n�0AIRi/D�������8��!Ǐ�15b4Q�0D�H�q�ߑsGĕ�bc��o24D#�-��hO�-`"��Pd8a��Y�+ͽeE�B䉏\�z�Ю�^TN`���J	�n6�=�S��M��Ϩy�X����t�dA���I�<qկ̌Y4t����9v-Љ:�GPX�T�_���!��v
&� ��_5� �k�.&D���T�����B#�i�&B&�Q"f�Ȉ��U�d貑��h\	e�����QT!!�� ����4k5 %L��.@�YK` �ϟ(�?E���	��Qe+�E�PQ���"�	��IA~�$+\��r��.�!Q�]��yҩVZ�
2��	�ԉJ@aA�(Ov(��'vܜ�C�RՃa�	(������l~��ӿ!��YZ7�փr ��+qق~Û����{��yW��P�y���;s���� I�hO<���_/-��C�AԈT���ii�Z}�	Y��hѷc@��Ճ�/Y�o4"�5!�O�O�-���ˤ AT��D�(�޼[2�O�!��ɋH� �\T떸���J�W/�B�Ix�T	HF�)G�v$X�n�}�\B�G�, ���L�>x��T�|dC���of�i�S�G*�C䉸*�j�q�kŕa�䁪6�%
�C�I,TŔA�d�U�Zkr5p��Y3#*B��5l�D���DF��v��9U�2B䉒^Π��6��1>-$Q���y����D{J~0�A�/��p3��$&\^�"�(�}�<9�$ԋn�6����)HB0q�@e�u�' ay�R�"���"�ْ��@�U����[H���EZ)ZN���b�(C�F-�ȓh�I�D�(E �Ad�߮<�j���Iq?O>��Q6��˙���e�f�<� �1Q"��A't��,b�ZM�I��ē�?����Ӻ#�"�:~�0pBA��-WK�ds ��R�<!&��9:T��@��*& �iD#�J�<Q�%��t�����#g�$�rW#F�<Q�痄	����7U�F�1��Z�'$�{��۷WV$y�c�	p#%��x��'��0�'-� Ⱥ��UI� 0y�l�ʓɬ�ڐ��|���P/ol80�ȓ2:�!0�)|(\��"�}�t\�ȓ\��8�G��|���oܺSB�q�>A�h<��Do��5V�Q�G�4�8Ѕē5;>�s��4X
.Y��"҈e��]���n�LF{�����'�`��n�%R���s�薙`p!�d;v�����FAG�H�8�'A�GўP��	�,���l̐S������϶�����(}�ǒ�_۲	��h��w��cd�@$@�B�+�F�j0�A�y��	��D�~b��?��}2D#ʧ �֬��D�A� �J�J�.T2��?����~b&Nʄi)����F�(`��dT�fyB��<�P�<�T>7�?5���14[�tC%%P� �h�@5lO�P��@�_ڎ�t ѣn'&|A���ē��=��0!g.�(��-��߻@�6���I8a8���R��+C��jՊ9��+C��y"�Јe\�9"L�+f|��")�+�0<a�鉙b:b��D%G�h���`�'bl�OH�=�}z��Z<I1/�R5���UCF�<�#d��0�!�@<`h���~��M�	ӓ�|�2�ŬzT�1
�I͆	z��?1	Ó�?��	]�>1�QO�32�a(�Mz(<�ߴ`��8�J�ȩ[E�wTd�ȓ{_�<���T�l��ddR>~��ȓD��B���#s.4�ч)��/����	5����gϑWBJ A�
�R��H�ȓ%���
Ү �as#�\)+��d�ȓU�~\��M��
��`�EE�)4��ЅȓmUȥR2
��p�CBm�0PÖԄ�Y6:a`�
�_>fY�P�Wx�*L���l��&lF�Cv(��̏�ff��F|b���B�2ˍ*t��MR�̈́�!�:C�	'htP�"�g�.���"S�C�)� �RlZ�60$�� ��U�>- �"O�9pB�yR���%/�6t�T��"O�kVIǴF&����G�Q��B"Or4�E�	�N_"@���>pqf��U"O�� ����a�π.+��̓�"O���U��'��j�E �n!���8�S�d�խv�H�8F(�rR���g�<��$*�S�OI�-saʪ1���d��/��|��{"��+�t2��2�S8$&5X�J�^ �C�Im����ۚj�4ъ�&]��f#<A��V=��V�t�L}�d��!j���C��'��O`���g��z��b5��q���8IW�'��6��m�q��LL�9� 	v!�0X��J�R)>����Tܓ��,�`.P�OG��pޜU �'=>EX@@/�)�'x�Y*�ߍ)�s�@�M{��=a�����E�!�z%j�Kt"���ĕ'�ē3����Q�Z�~����:w4s��S1�!�䖛7.:�d�l^J�*b��OW!��;F�RL�&f��=P2�85#��TB�����y2����=�f���JF��Id3M�@��'s1Ob�#!�%�f����0|e�1�|�)�ӘP���"P�vH��FS~B��=s*�	�NG9	�lx2b'U?"�:B�� ����F	ŉ9qMq��SVtB�	K3�P�!�A R���1��ԴH�*C�	�i¸)�$�!V�ҡ����
��3b^��&�D�	F��w��nblC�	�D{�hq�%Q3���cG�G��Op��^ܓ��'����c��!��",H�6�э�>Q������ȥǅ.7D3��
O�!�'!�2�C�'�,`dE��)	ў�ቤ;��}�t(�;��Eۢ�H,��B�ɰhF�LY�Ê�i�ԥ�ь�,�^B�I���s@��J�X�@��R+ ���5�d��i0��	M I iCE��&���>�e$�NYƁ�孇�Dk�)���z�'�ў�$��q�"V�!��HĠ���� �Nr,��	O�7�9�ȓB��j��ֶ(B�G�4dy��ȓX�� I`LՌqCPP��#�+�$C��
6[�)���;n����kL�Z'rB�I���qW.I�IG���,�zHb���ɴT��9)W-�U�����k�{֓Oޢ=�}�3/�",����R����L�
ԫRx�<��톇r�̨�q�K;r�F�k6k�t�<6�O bp���A`�B]��F�q�<�R R2:�Ҩ�4�y�MI�K�a�<	b�	�`)3��H��Ybe[T؟���",��#jе<�b��̙�N7�\�Op��ϩr���b��&u�V�h��Jy=a}"�&?�@�Vv�a!>͖A���<�6.�!-�hq�3�K�;�d�o�O�<	�ל;T�P�A��V"�0�J�<���L�,�b��ԡǞ/p��)j�<Y@�޾�s�_�*���pĆ|�<�u�E*�a���bŞD@f`�y�<Aǧ�0Zt%�D�Ďb��ܣ�MM�<q�P� )�a�poYO�ԁ���
K�<14�F�:�)��F��NP�Q�G�<`/�w�>!r�-b���:��W[�<QaB�!]�,���p]���TQ�<1�Ƙ�:4 ��D"�l"�К��K�<��b�>�>4)6�W�N��:`�H�<�"�_8�+pϚ�!.�A86Di�<� �u���1+fjx��,n���D"O��%�(��&n�m����"O��tB�k���NK�Ec�%Z"O< �J�OV��A�O:(|�(�p"O�$B1��*169�T��me�
6"OZ�h�a� $�֩X:
A�S"O���ń ˠ�@�h�)*r�"O�4�"J2\� �`��'�h�6"OZq�g*���XWOV?�*�5"O����*	;�Z�`a�^y�ȑR"O����@)ܐ�߆&^t���"O�ᒦ�Ø�B|�,�-�H���"O�Y�"�'�@h�6��	j���8�"ORa��BTm׆���<[��@hU"O��qaN�� ܩF��u�����"O�0b�W"k>BQ��V�M�5�b"O�0���M�x&�ly1�ǃP�q��"O��"5$�t�3���F(aC"O4(`�ʀ�U�
}+�)	�/c`Y�R"O��� =�ʝ���%_G�e�"O,X��	��T�ʓ�E�y$��"Oj ���I�30<�
�F[�!5QS�cy*	Q��GZ.�T3��E!!e4�	���0�t��DEֈ{ѣի��B�z+P�1�AH1���j�kt�BB�	;��P�g�.p&ḷ�hʂktC�I�L)9��Y=Y B(�b�H�J��B�ɚT���E\���i�n]��B䉫lc��k÷,8�!#��8pd�B䉒>���q�@K-�nŰ�)
��`B�I/_��R�څ<�J��`!RâB�	2i�v}Zì]:w����P�о'!�B�({���������O�hB�I8ň��G�Z�yˇ`QS*jB�Im���A�&��1���� &6C䉳p��EsCL�9����ԍL5w�C�ɸkl�Ua$fӋCD)QP�	9V�B�	�Ut�b�(��~fM����\��B��:��Q"AgĎj����f�!J��B�I�p� �K���Y}����/O#��C�ɩ	��(��kG2HC�Y��獒-�C�I%h��13G���a��(�AЊC�	1k�ܥ )�)2c�� �)?fC�	�rA1�0Cx���cBW�hC�	1Pڢݡb,@�E�j�05�-�pC�I6_�=x#f�[h���G
�C�TC�I�q�Y�P�ů�b}�2��J�4C�-(�> Qf��Wz�!���B�	$
��1��˂_��Y­ٟn��C�	�~A>EG ^�t	�T�Ը�,C�ɭ9������_����SnӛKG,C�I!o��21�*	�#l�Oa�B��?�6T8v�Ο]֬��ʎ���B䉈%\���f�S�92$ʑ��B��2-��k�L���p�DF TZ�B�	2_4h��M�sp�mA3�S�y5�B�	+��	 f*R/�`��o�B�ɭh����EI�>v�j��R�R�*B��=AѶ KU���S<PA�SO�$G&B�I�y@4�����<�hT����C�I:_RH 豹��b�[!{��5�s��<'~ȵ�������␈�(oܠ�����G/�C�	$n^�0�%�2sĬ C1b��fEy�ŏpY��Ob�}��)���
�_���B��:P
R��?7D h�!�-E��5�t����o��$�hS?$��{
� BI�$�[�~��c��Ŭ�°z �'oД�Ń��S����w!����BQ�*�T!�e�2^��B�	�l�����Y�E0$��,u�Hb�Y��\0� �Y�;G� r��Шc���r	չT�JB�I�2��\s�
����MKvL�3<c*(Q�,� �~�O�HD��O0��a�*9�b@)!�B2hFᰲ"O�1ӃZ����&�4{e@T��iy����+Vت���	-��F�B���Б��IL���$��9�6)1�`�4�?	T(Ӏn�^c5�E#i��x�Y�<�j�#ٌ��!�Q���`v�OV�Ϧ�ْ������yH�L���$��"�'�Pd"O|��E�9O}�H��$��
�:! �"Oze)��ˉù0�ˑ�Dl3�"O֍`��Ϭ�Ty�ϗ59>Ų�"O���� 44W�5�#��c�МB�"O�(�)X�_T�Q�B/�Q��"O�=�%�B#px��qT�M$"lq��"O��M�<5_��W�/�(��"O�]q��]"6�����Zj6�z@n��'�qOr9(��Y���Ƌ:6�����O<O�BY��-W�l��O��F��'0Lx����>���M��f����ICF:$��hX�x�B�ԫ\��͘��J39�$C&l��.�B����;ʓ_�����J2;�"S6Lt��p�M'gvH��ˏ�%)̩P�9\O|��)����dA�*�*H� ��w� �2�_R�	U� )��L>/�<�b�E�O�h	���@��#�����@�Ѝ{�-	�x+H��ᓸldyV�|T@H	��á���eQ�m�Iu�8A!?�3�	5~\ӢaͶ7_2,Ǐ ('@Н��'�I�#�Q>7m��4	t|����U��8U�8��]�-�а�0�s~�[ۓAV|
1MI�Pf��w �2�X�D�&Ԟ|�?�T��L4��C�A0c����j�=�1�D(�X�R�ϙK����m-lO��C	8}"ȋ2���Sq��-��@�6.���
**<p��5=)`)Q��Y�~B��'<R���kh>�[SL[
Y���/I#[��bӮ+��K�M'4�,�u�tه@W2y��|��B�*h�x�B�!Hd�׫ʔO#0���@1O@���ʞ�N�,����ZUA��OXѻ�IU�W�pY�'aj�rq�T!@��Л!Mا0͖���ɇ4�@=Z䋈>ޒUJ�̉I�x�I�?�J�� T�l	�݈��Q
ƨ\�'�=��c_�B/ ���8U`��m9��$�)���ҜS��l���;#��0��ڊc�(�1�')��B�ŞV��Y���)�H���z��q�^��Ԉz �D�Y#��"(U��Q��o��P�w��p��G���K��38 A�U��X�$M�-S�l�q�
�yp�x�$�Zŋ�!/��� aH��|���S�P�h��+�9�Oφ~���+ �i	`m�hP�|!7NV���OD�0���sI�Ua�'̦aQ�����	x�A�:ʶ���9'����PjA���ÌۊV��K�L,��9��d��1�@k�J�3�*B��Ɉ{�mz�O���\�;N �í��[}6�`�].�eȠIʢ[	��p�S	 �a�5$���������>	wg��$�zP���I��������*���I�
	�q�e>q��\9'�A�!�b`��`_�Z]@�[�Լ+ G--fjx�c�L�Y�N���~<! �,1��e��T5�j飦���K��%k3�[�"�FM�1��n��T.11��m*��e��LR�u�Τn��6LDA�W� Sy��,�)w���d��_#D�O��P��)i�\ȏN�Ai4�Ɠ?^��V��s����H�E�d �#�(j�RGz"ľ;O|ˢd.f�Yr'��p<�ulK@��a&!�=HY(�O�+V�|��c"���p��G�u�6�R���88.�\!	�7���MN)Үmi�A��%�hҦ	D�@��ao͑8���rq-�o�J�$Z?1���1_k��RC��~��a+��9D��t�N�;�J�!�*�*w��2�d�H���U�|C%L	����9Q�wg� �q)T*'�漡�d	���'����C$�0<��Y�3jJ�iN,��iX�9E1OL$�Zwo�">�pDS;DA��3G�1;n�;��_W�<�� ��o��P�BFy��,+r�[v�<A���A0��ؕ�F�eڦ��q)�E�h�~P	Ǔ��eb�I��';����"%j"���z�<1j6B�+I���is�@�ɋ��"e&�C��5g>`��Þ-y�:9�5HϣV��K~����y"m�p���Q���@ �Js��-�yr�,z���3q�ܒ;m��.���8&|�R���� �)�A�G;Q"U��%�?D0��"OV� "C��ĵ8$���,4:%�F�����T;Ód�p�]�t?�Ų�D�i����|���'&�y1��k��QI�"�B�	�������"�x���~	d��D��)@➀*F�͠(`�,!�JËI��`$$D�(��M�>�)`�� �/f��qH�Bܓ3ʎ�(���x"㉏<X����K�,�uϑ��Px�G�]��P'� �d�8��9g^��`Xt3ae�K��u����yV���%�0<i�,
�ԓ�
-}��d��:6�L��E���V>�y��Ѡlo$(�Fփ,��Xȉ2��D��Q��I0���)�'^ �"5�G�	�2e�c� �`,�ȓz �b���Ѹb�i
 ��gA"}Re��0����yR#!o�Xf��'�����Z��xr�� j�\��F�]�Z�A&����`�aͦ=k>������(Y3�ӿX ؍���l����B���b`����4L�@f��?��A��
ӫ0�<C�	=��!�N�o�D%I��P'6
�Q���2��Mhҧ�J�[OT5RwX��2�M!��$�"O8��@%� #A����)�,���I<$��#�9�3才�=B��S�Eb�̜ 4��C�	u����P�}7`�@c� အ�aљ�����ap&ϒ�7%�w�0J���d% mN�)J>�M�A�t�U�M�,��`���p�<qF%R�Zj�p��RT�\��kZU�<�p�K+$4�2WlL0�@}����H�<��@6	�-���a��A�'���p<I��	'��'�f�Q$�V��T#U�^�s� �Q�'*0�7�C� R����׉\q:�O�0o������"�x���{I�Y�P��?@����"O�`�aFW�5ވ+֍�v2^�9���s9J�!�t�ݣDZ�S�530k�03m8؆�v������m�"�('�խPsa�vD%)�B�I+T�^�;�̝iOna��G z�����5o�Pc�{҂�(E�9Q��D�K�y��Ύ��y���\Dt)Xp%jKW2Q��KL-���
�+��p��{�������⑏ևH7��0��w!�$#��ݘ�����*�����ڀ��
G�p��䎰>�-��`F�U/t�y1��e!�d�՜�����<�hx���� 1!��3\0�ƍǇi��I��+w�!��7��RgŠy2$58��d&!�$�sr}v�ۗvD"��d��-E~前n]���
�c���	�X] ���C�	���c�
D����$G��*�A0�K�C����<Q����S���$�AA�J��?q�L,y�jŁ��ڔJ�`,���w�'=JmC��-z�l�����R���T�#Z�����K�Іȓ8K�4(�.�p�-��,���E��Dς�fhH�@�|�$=��������NLB���Fъ2Ѱ�Z�NX��y���#�:)Zȕ�)|h�ӓh�_	���#v�D��bg�>��tȥ�I#�V��@Mvz�ш��L
�z��dև1S0���%H&W @!�l��5�B|&�ã�z��t�ԣ��rD�&9J�ER�@�����1�9�(O�k���%?@�Qbm����OX:`c�H�#L�a#Ǩ�nH��'�:���+�6פ�"��`�i@�Sz�fA1����)��AǑ�v�����b�2)�8B�%D�hrҁ[�#��G���zS`�f%��qЯG�	{�����'��Ҵ"ͽR�|e��)J/~wV!I�^��j �@��؂�
eE� ���NjG�c"O~����`}���ǒ ^j%H'�ɼ^�><Ss��}�	sΘ6"���L7g��C�	 7�X��"����M��,[�x��C�	�o��a�v'��:ĢL���Yl��C�)� 
#�/D+����DE��y��8�"O�TKgᖱV$iC$�={U����"O��E��6�HYPcC��o ΍��"O� ���Ns>$��bևJ(]""Ol��2I�%0�Ԭ�AJ/Y�P�"O��k�?&�Z�P�(�TuR"O0��KW�p���&hQ)KP1J�"O<<*%p�Z��RGٕ,��Œ�"O�0a&Ð�DE扢��=IxD��"O��'bȈ��I����1�95"O�U8�h��K�� 1 �_&t��9K�"On5�Ȋ�MQHt#��[e��"O�� Z�V�T�11AդV6B�c�"O�%��݀��4!��\�*j��"O���cI�2���5OΩz!P)�"O�Ȱ ��<�۱R/���"O��f`Y�]��m�W���\U"O�K# Z�`=� e�۬8�L�XR"O�+ŗx%��qr��e��Q�P"O���T��)h�<�b�̭R���yҋ�;@i*�Q�Ǿt�Tp9&��y2�F�~��ģQ;����M�y��şva�Q��D�^*X1� ݨ�y�j��Y���`�ʀJH����#���y�Jוe:n�3	�)EJ|ؘ��Ж�yr��=�V�#@̌>�RUc"�ۅ�yR(S�|H��c�6���æ+�<�yb!���h���%p	��%�y��0'��$+��`%bUNS��y� �/����p,CX�����@&�yr��.\O�q#ޞW�bT&���y��B+�f(�\xR<љT,��yR�WФS���;F��ɱdm�y�@��;b���cR�!˜�@!�y�F�8[�j59&.@$mF �)L��yR�"r:�Ț���&H�A�����y��$yt��c�C� E)U��y��0*������:��YBu�P��y��3��c��c��D����yҦ�O��p`Pk
Rpl$��`��y��*m�R �lP�Z��1�W�I��y"��9�5i��)V�A�"ۊ�yR�O���5P��[��� 4�y�+�;xd�� e�ȷ$t�-�gA^6�y��L&FQJ�����$�\m!���y�*ąU`	׮�/A��9��_��y���>+�ε�s�\?)�i��n�/�yb�zh`��!V<��Η�y�I�"��!!G&_�!iGd�y�@�cr�1@�W�ȵJ�� �yO�o���Id��+T�(Pf�	�yR�]ؠ����'�Ȉ2ukF��y�,��f����n�"ERD�t��%�yY�lM`�)���2"��J�-�y҇�'Cδ���1-��0Yc�[>�y�O'��Q���IH�z��P7�y� �0[�e�G�Ή8J�eٴBϩ�yR�~i�� HpX���D!2ՅȓA��HJeƀ/{{�Ire�!\S���ȓ0i\I#D��4:m.����X��|Ņ�f�&y��U�L��87�c��	�ȓokAaF�G=|�*�e#���ȓb�B��O�k�D�zr%!��x�ȓs^�����O����/E�
>��Gxr�����E�� Ҡ�&6c� ����,A7�,��"O�z����\[���H�v��(�+�����|"����V>��L�1���f��-��%=D�Ȑ7�ֵ+�i�SE�)cCixӂ͂6 �h|�\2��4@�2dZL9���ƚ'>b���	#]_t� �Ʈ\B�
�2�.�R/�g�r���)�yr��f�Ĥk��� P�t�r���$��'�� �� Q�qG�D��;�BMpEc\6evD�"�ǭ�yR���{��Bᮙ�]P�|iB��9.d��iޢ��q��>�
3d9�a�@@���r��/8�,��.�j�*4
�Y�B-��I�T���m��U�P	�K�*f��{�ɝ�x����,[H���@�H���=�5�	�f��'�O�#�M��\�x�� Ttb�	��"OޅB�(�k ��X�`؎@�q{��D�5lL2�+�1�t�����M"�����5E�d�ȓ;"���D
͛�F�c�̈2a�f��ȓ�%�`���P���ͦ�����5'�b�65��%�w��Q��d��Ci�&
��q"ā5Lx���A�6u26�ٳH��H���#�0-��,`~���$ch�t��ܖaB�Y��@M�pC� "j�5�
�H����V�Z�,�Z���[n]2���K"p��T�B%�8v W��|��ȓ�U[��g��Њփ.%����$�u���	&r�v���*Lr�x��Kr r׮�� �p��앯<�zY�ȓ�8�rW'	�D�M���ݧ 6�d��v��@�����yX�K�]K����L� �7(
�h���C�*ɘд|��9��Mrcč�3�uжG	�3H}�����瘗m|$mP�IE�3�V5��D����Fqv G�B/e%�D�ȓ��,��H�f ���*"��X��B��a�0\�uZ�)طdO�P��=Q��ӂ������4�Hb�ϛ1G�|}�VD9U!�䟔6�E;��C+2X�ȷ�P1 `�2��aX>��dٮ^�>|a!CL���6d�='�џ��EE�2>,�s������AvL�a�
e���Q�!��^��a�!G�:mڲFK� � �'��(�P��L�dҵ߄@N��i.O6�B	V,y)N�d�Š�/_�.z",γIBDؐ��4q��@2���yЍ��%ڋ�B�	� {��!���I�I�2@S��B���I4�(I���5 �$zţ���As	n��I̻3��&���;CLʨ�̫�/=�O։-9R� ��;G����D�6�&���< �l���	�)WP<I�OҙG�N�CPLF{�)�%1�D��I�HEa��VȞ�p�� `�?ADeMJ�B	CR�=�	��Y���	�9?С������܆m|����C�y�qaN	��iDzb�� j����Ǚ�tM��-���d�oj(��C��ē9��xd+Clczp㖠6 ��q)2+з��X",K��.��Yy�+Q�	�a}BL�5�n��i҂	�h�E���_���'�F��/S������ю9�"Q
���k���b�;�R���֘,%���3��̩vOP�8�Mώ�pa��3JiJ2 +���ШpA�n��4�� �T)�qK���d�2P��M�A�9lT��� Gۨ_������n8�T�Ãl��'�pH�i��u��;��T����i �@�"��j�@��@���ꊚ�dxMa�'�4\��fX�yBE΂�@Ժ�iӓ,�4�
7�ݠj]�<J�A���#q�˛HT�
���g�:U�q��8-�����'���A���� 2q�H�+��{2HZ�	�I�o�I�IC�D��I1pP?�ER��J�!�Ԝ���b��9D��b�Hԋ.�a� ��	jW�	p�9�	kS�X���j�OF���oS����'�	EN���'����֝��t�$�;CVȊ��Z0��'*`�E�,O~�ӱ�u��;�.5.��×"O��
��w�&��G�H �DP�7"Oh�!֊�-{��I	��ov����"Ol<q�$��;��8�ib��(�"O� �1@�$+�D��1県)A���"Or[���@���(4�U9e:D"O$
���'�����@(BL���"O��y�!"@�h��e�I�D�j"O�,9�j�"���qC�U� Q�$"O�@����@6d�(-x�;"O�`tCX�%Z����n� jP"O> �'?+J������i�X��p"Of���92d8!m�*10P"OdhSb(�-h��{6MY����"O��{ /���d�Z\y_~���@��'�܉�@�%�3�$�28n���É?NE�q�-���D�5j���OܻS0�1 @;=���au /�����W.9㓢R/mM䩢�F�@�axb�Y��tu[rUe��I8��UN� \R�1�!��7!��rg�a�A�X�:�;���u4�	>F�B]��F� =��S�O~Z���u����(Bc���[	�'��T�ǻ���(0kT��pA^p���cܰdc��?�D� 7x&�3"�r!��X�|�*]Y'�GAcj\�6�F*q��Y�� �s�v` �+)d�pF3A��P 7	�쥇�	�Y�9����9Kz���5"��ZG~Ի �Y$UYr��k���X'�A@�H��ǉ@�����'�<��ϒ�\y�O>�`��wB�jB��Exa���4D��a�:ߢ8��ȃ��@�5F,g�3�ȹ���M�g�kh��HFn,8��6.�3�l\�4�zL�1%��\��bG'-O6���V:�s��&J]"Gƈ~�,��E��'a���I���Q8��|
<h	�A��E[��r���y����d�]3c�e/�P�h��y��S	T�
a
��_Z�9b�2�y2�*B��!�
�[{\��Y�yr���@�v�#Ê��R��Ѓ�e^�y2� �1t�$"3�R+ �)�����y@�r�,�����.`HRVgB�y2��"M�� 	�PH�9��@��y"JMF(���A��X���L�)�y��'M�pCc�'U"J�����y�%�	?���q��QV�,�*�C���y"A�%irX	�a� J��!0�����yR".P������@v�z��Y��ybQ l�b!K6�5U�^�6Ǚ��y�c��H���P��th���Ĕ��y��ʘ~�>\���s���7�ì�y�C-3d��xҍZ0\?>� /��y�e�-F�M���"i�t�Ǥ;�yRƸ���Z1cW 8�C�Ã��y�jگhH��G&�$|62A�L���䞙A����ۓOhv`�R7~����׌�,o�u��I�X>�ôI�i�[R��t0(+�i�1B�bB�'z�l!��0v?|���G�o�و�|�p�C����V!RS�Ř<�ޔjՍ�-����"Oa
��E�T/Pz�Ƥ=��<�`F��R]J�Uġ%��S��? BPP��Ib៻,�X��k�U�<���0��M C!�1,���ˆ��k?�f��E�IY�O<LO0�괮	]��S��Ċi�ʵ��')��z��)I�0��V�+7�
�*�8K�@�G�H`�<�3�OSҼ�E���1^�S7Va�'j	���JTشF�doёg�
\j�K�*@*�E���y2��T��XB�EL�������;3Üqկ'aW���L�"~�ɜ
%`p	`g�86N�9�%�$5��B�I�'�:1dC�P$z�pV	F.�T�I �ʜ�ĲK1az���;�h�3���<@[R� ��>��$@�.��bGq�`�R!H4`��� �� "O� �*��R�rD��"�,� p�t�3���D�S U�\tjI L��]K��U�qE�C�I�1���!a�*��%�㏑�`B�B��U'�(ԍ˷_�j@��O�XʢB�	�p��,ic?BPT���޲B�	~A`�cU�Zjb9���#<�nB�3h��I(q�@�8�hE��7M�VB�	Va����#����%��
��C�I�4@X0�Fj�
G�M�"��B�ɖ9��AbT�z8v0B5���B�I4JCH���KJ�$�\��#L3ǘB�	�\����X7QA5��+Ȯ.�JB�	�D��Ô��;�T�A�H�K,B�I�l/"�� eiD�U�/4TZC�I�]R�C����k[R%��/�4�B��=/$�y�R�M�l�C��wQ�B䉀i�*� t?Oܨ4�$If�C�	n��cb�� P.I��_$Q�C�F���%��}Mɪ��]w��C�IfдQ���߄-'|��� 'zB��+91v����.{'�9�#��dPB�I�o���b銁,�ᣖ
� B��,��׭\",`-zAGK�Y�.C��R��w W�t�}0D�K5�4C�2� +'�� g�.�9�(F�:C�	�z�q�a?F(15�ǋ2�C䉴	`@Y�2-��ixi2�BE.Z��C�.F��˥� �m?�4�Rm�s�nC�,Uh(�&�=+�А��@�S[�B�+IR��K�s8�<����e��">	թK�3h����@� Q�W�<�3��:bPP`ې:J��k�o�P�<����W�
�� ���ٛv�UM�<���
9����3�أ%ʇN�<y�����(������x;+�K�<a�m��F��-�6B�e�.i#�"_b�<1�H�4~���i i��V��s]�<YC��r���yf%��u{��TD�HO�"}Z]w���I�:|�F�a�,�6֎Y"��T���'�
d3����#_�(�@c�ϕ���<�G����'��8�I��O�j��O�8��R��`2� gOU

څ��'\S�IE�{�PT�O�>=�K�����s 2��%˒�ڃ9a��Ñ+ٚ;`ҧ����с߁y�L�)��֪{���������x�I7�v\�q�,g��R'E��`�K���'�b���qO�V��)2�Q3g����BK"#5�X�<��b���<�� �L�=��m��~�8����G�<y7�[�.@ q@�G؄$��a����@�<A��I4`��m a$Ή"�~Ѩ�M�Q�<��H��@0 �ӏZ<y20ݸV��M�<A���={q�a�kU:fd�`pL�LX��O�{��D9>�)�MF����"O�u��c�mR���-؏���&"O�����KiTu�B�J�G�r��"Ol� Q�
hA(�K��e�"O�a%�8~/�(�iM��%���y"�"i�tu�u2� 	ʡ���yrʐ�6��A�Am�<��pP��y�B�]t�)P�;zt p��6�y��~���JA���ƕ1"㗽�yi.FzB��T�׸'�V�dW��y��R>�z|�Ӥ����lK�'�(�y�!׳=��(�#l
� Y�ԧ�y�F�d6�;E�~=6�* Ŝ��y���d��!*�N� %(�T�����yB@\J����Gظ-=�)�m��y
� :̀ ��>	W���p�I� �Ra�"O��s.Y!�;���i�V\�q"O�]����XG��Y��@� �>���"O���҆*�Bt벅ӫs&�)1"Op��䆊�+	��qU%/s�pa"O-s���3\T� jV Hq�E"Oʰ�c����n��ň!ϩ,�!��N�~&0Yyg/	�'��tc���9z�!����eŅ=����n�!��%�*ya4/ßR��(%@�Xg!�Č��j!Ҧ�3dh�A���'!�$N	">T94��q�^$C"˜�9
!�D�B���/� H�dUD���!�d +�hq��+�����B��`�!��+]Q�'�.'~�)��()�!�Ĕ0���y@f�#��`�g$�2u!���2�|,R�V�r1  �G&Q9Id!��]�Z�`�!U�mH`Hs ,߃k'!��̈ |�Q��e z;��.T��@"O�0�f�ψ)�F˧c]�`/�Ap"O�D�e��/y���C��X��Jq"O\���#�X�ɱ�b�%o-)��"O���� \�><��a�Q�ɢ6"O�P�TC�(1��T�w���P"O��(1� ���cǢ)�(E{v"Ot5cU&���y
E!ԉr�nHh�"Ot1P2+�O��!�T�0��s�"Oح����8���d����G"O� ��CD$�"�$ ~԰���"O��.ӷfY$���6�ʀ"O�@R2 M2������5Bb䍸6"O�d/ o���R�CU@T��"O~ͳ��Ơ���(�*�VOPر""O����M&` � S� ;~DH�"OB�"�-J	@E��@����M�"O��X���w����'��y=����"OrI�鏆i3�uJ���� "O(hK���8E�E�"��! -� "O�:t�M,
� Պg��n��uj�"O.X!&��\�8���+?��(�"O�y1&��)/h�c"�F)�P��"OV	�ӄV'\��lc�J�,��=�Q"OF�ͧvz��p�$|�t"OҜ�C�H3+�NLR-I%E|�U��"O8�2�V,q�� 3��ܘQ�d��B"O�q�a��K[ ���]KY���"OH<�c��$�!��jG���u"O�x�Ɂ`�HYîזX*Xs"O�Eɤ��S]�A��QY���T"OJ�"G�,'2\ʂE��m�v�у"O�]�KK�?���sʇ>iJ �B�"Oؙ�c��&&LzQj�+7�AQB"O@���hB6g���C�ԉG��u�e"Od�vH��i�~L���I��.|�"OtX�! \�T}z1�۰}�Z���"O�	{�M�7�(��NI �L(S"O�:Q��i�M�d-*(X S�"ON��!Էj�(r1L�HR
�"O��`�g��� Fj� (��qa�"O^8 �eƇ��5�[<I��x�U"O`��C�8G��J�iX�w�<���"O*Y4넲�&\!��(_�v]Bf"Ot9���Y�)�Ft�6�	�`y\�g"O�h`@`��~�&��4v�IK�"O� ԭ�c�C�d�Pe/ �}�p"Oe؅���H%Xx��f߁J��Y�7"O� ���tA*��B�.�b�"OF��g�3� yi��Z�y���Yq"O�H�1�T�vr��@"��nK�"O��P!�X�G܍��;>�&p("O���S ��K�Zd�� �>��"Ol԰��O�U��bF�>���P""O��բ��N�
�[��� w��B"O0��� 8?��q&�{$��"OF8�Ŋ\��,tHV��H�t+1"O�i�S��-N3��R�c�⥌��y���"ٚ��ւ|_N1󀭌��y�,ūxi�Ǡ�>s����`O��y�'��M�b��#ɭh�
Q�[:�y��[+L�^� G�G�8(i�n޲�PyBo	îı�#��	vR$Ұ��U�<��Hʴ#q<	G� (������DN�<Q��37��xa �
(
{��!eM�F�<�e
^�^4����b�$1[�	�1
�H�<�#�`�KJ-L��5�� 5�B�+����� ю���F�g�dB�I�h����$�����	)��B���`KB���j�_	H0*"O�#�́FȀ�B�a�"����"O��C�R
ng��o�Al=c�"Oq�v�ʛ1�"m9D�J�$[��R"O�\3�hoX%KM�8<Z@�5"O��z�F_Q\I�a�n0�x�"OV ۅKR0u|�r1-��r���"O�5���R̄��'��]�~�# "OjŢ���IEH|8�͂:�Ή�"O(�4�&i��8���A�z8s�"O��:����8����ք� Q����"OD���C�5qh�D*�c&R{���t"O8��T��Nƭ�2��qҠ= �"Oe["F� >���FO�.*v�`!"O�eB��ŭ5�5;��_7k), ��"O��3�� %�:�
���+���j�"O2��g<(*�{�Μ�Ba�݈�"O�T���/ό᫰�C�.=��7"Ob�('���B!ԑ{EbɥuW��+C"O���2i�
���ɶ��)c��yW"O2�	�/߼u]f���*��^����"O���K�H��!C�K�%y,�"C"O@U�V�]D=�li�H!F8H"T"Od 	��	w��W�	8�Xc�"O�Id� ';�\:�)�5$���"OhAw��v|l��3�݂J�`��"O@��W�;6��sS��s%"O*E�̋8R�������
l�xh��"OTݳ�Y'Aټp�Ƌ�<(�Փ�"O�Ѩ�3%OZ��p�@�=Z��"OP�@靅��� ��0KX�i��"O,S�� ��T���HMT��"O�� ���+De�vNU2@BipW"Ov���R�.��@�#L�&RZ�@"O�S����p�#�k��h�1"O�4�s�ˇ�jL34�)o�r�z`"O25j��W�9"d�)�#N�Y�f\X"Ol��KB�1�8`��ƀ~3$�;W"O�d�w�ru˶$S�a�6�3�"OP���$V5i��%87	ɭ}��̂3"O�eʶ�-3�xxrbK�l���K�"O� Dm��N�	x.��C2��9"Op�[�K.4�>�p�i���"O�(��,��z�j�p@���z�H��"Ob���n�0TM�@�Qu¸1t"O����aC�'�h��p훊Qc+T"O�X�GCǐ,���ᆢ�8^F]K�"O6�q��Q?��%��@^5mL
"�"O
 PA�[<@�eE����C"O�h���._�.��<ĝ��"OB�j�D��eQ�u3�o��]��"O	F�$_��i�!�[>P� "O��;�kV�z\�1N�/>a�x��"O:	3�zP��8�M�,X�x�@"O��6f����	u�V�M>�Q�"O���ҒE�h8�O�&*A�8�&"O���rg�(�JQP�OR	6� �1"O�$A�+�<نP�F�]�,�R"O�1����C� c��J���"O���.J�g�(� 0���~�ԝ1F"O,�##
��	�h0{�ā.�ȭ�"O�0:�V'�&��CJ�{�|�q"O⸉�i��w_�}3e��*���XT"OZ�yE��!)Q�8��O?_�0<�r"O�1;�g[�cA~`!w色e�j�Y`"O�QI��ӥ\MRL	��A:�R�$�y�"�/�Lڂ`զ\O��K��2�yB�!I��ɳ�B)RZ~�`� ���yҤ^@��MJAZ1E��yk�(�/�y��@�L��A��t��@��y���<!��=)��/�n̰5胯�y��Nx}l���T%~��t���yB��.�Jh+��t��K�CB��yRE�?��ac@GJ�(��Xc����y2,ݥ6d9��
�7m�肶OT �ybk�<���2^L�x#!-��y�מC�z1��ң
^�=k���"�y��+p(��_�}��;���yb�� x9
�#�D�K L ����y2j˻<���	�[��P�Cꐶ�y�*U�l`�������:1B�y�C���@8a�*j|I1�y+�jМ@��W$�|R �[:�y�!��3�p�����d	��c�
P!�y�W�Y 3�O�PqC�I���y�B�y_�d��Q�|�b�� ��y�&�&W��"v#�s|������yr'6���M�1s�J����y�aS.�Peօ�5^q��S#W:�y�ᄁ1^�53�o��X+����&�yB�Eb�tC�(S�K(\@0cm�y���c."����X�B����G:�y�	A�f� @"�&^8��ł�b�yr�K����j��Q7�.���'���y�ǁ��>�ȗm�6vP�EY��yBG�^����#��%\ �թE��yr��2=\t�i�X�mP�ɧ��yR��$|�.�a�!��.�����y�U;�9�c�	�,Ȳ�"�y�̟�A���h�����p�E��yR�G� P  ��   �  `  �  L   �-  �:  �H  �V  Vd  .q  �}  �  �  v�  z�  �  :�  ��  ҽ  �  w�  �  ��  �  h�  ��  �  b�  ��  � '
 � � � d% �/ 7 �= G �M U O[ �a �d  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf"O�Ya��=!l���Ɔ�b�V��!"O�!)��Y�fx���eE\z0	J�"O>��pg�0Z�2=�C�A�Hy�"Ob\B��;h�`��Ɇ*���S"O�h�T�ÕZ(jܫ� ��+�Ƚa""O�A���I�{"��qReM.v�\�J"O�I��cR�G�Fm+De����(�"Ov�M�{�Ҵ�U���F�T���'�Ib�R�HV]YT�i2��"O�Gc!��̕��ݨ���i�	�!E� H���O�6��O� ��S����Қw(��֙5�mS!���~,!���lib9�3�D$"wx`��b1�ơm~2��`G}bƅ�>��%g��	=^%3@�	*�0>�N>�ԧ��N?���Ý	K��`���^�<�׉N�d�d����:+�U��^�<�5
K76d�Ve��X��8�e��]�<�b�іQ�d��UL&O㪄;���C�<��N��7D���K��Z���H�G�E�<�a@T�S�M�C��`���"�C�<��+��6
��0�G� ?����g�<9�A^�t2�=3wG܌	OH�<�$�^ ��Y���M�w�$��Ҡ�L�<���ѵ.g�]5�	��Z��U�d�<� �h�-�1*�"�ѵk��E+�\��"O��q�M�{� I)�	Φt ���#"Op����G�(�t��5�2Q�z���"Ou�b��+Aj�"W�SL��CF"O��u��5dPxW�-��Qf"O��s�];(��q�#di��2�'��I�*�^@�O�NU R���0bP��p?��Ti:�B��Il�̑C�'�a�d"�1���0,I�{��u2�F7�y�ٻe�Ԉrf(�d`�i��HO�u��SP(ę���+b$��6Fl=�C�I:Y>�a�A�3=đ��oD]C�ɜ�h���ɓ�ڈ �e�:�#>��R������2!R�����V�w�����'�Y�<9G	���h(����g�^�ieT?���O��}}R�?Vy�l�ݚ/���`
�y"bQ2�:tP��R55\J������UX��2��$1sT="�$�U<�t$;D�����]:RZ򱙖�֯w� �x��:D��(�jH�cP�s@8���7D�J5�S�3��QU�ϔ؍!��E�<�/.�J�:�Jа7o�Iye�[�<���]~��Ɛ,axd�� �R�<� ��H�X�M?$_���2��b�<�"��&��퓵o8c��@��'ED�<�f�.>�<	�W3U�|�3�T|�<Av�B�l��H+��T3Yҹ�BHz�<٥A� F�j�RtoO�/ȆD���P�<y�G%8Ŷ!ic,]))�r�Qc�Tg�<IV�R&��VF(0+�]�p��e�<���ӰrW���J�oླྀ�jRl�<	�AM�o^0�!G0O�d(�`�f�<��`�/`g� o�<��@�g�a�<�f�հE5452煂�t#h�ad��b�<��6K��Q��A؇B�,���SU�<I���Si��1 �	X�`�9îQ\�<9E�,-��sB��;��q�$�p�<i7�!q8��R��>_����&��p�<	��L����	�3�y6Fj�<Y��Ϧ�T=�d�S��|p�Ye�<Y�ɮz��}C��V"Pd(X��`�<�bd7]؞�!Х��c3V`@2g�S�<�ʹ%��Ձ&ݦ?��P�n�R�<��#ӇT�j��-"���@`NO�<aŭH/R�	��W�B�3��R�<�'� *��ʇ
� X�䍻怈O�<�!
ַXM���HU1=ɨ%s��D�<��F��C<�͚�)�\����
C�<)W��#[0�T9𡄤B�L�B��~�<)���3�x����R�v�B�c�t�<����3�r�J���[Φ�[��Ps�<$$�h�x�Q��p��P#���l�<iҎ�
�bh��V�jm��a�g�<�ńS `�LI�b��!� jr�}�<ya�MI(��T�ȯK�,г	�w�<Y��ȿs������L��e�l�<��W< "�9fD['s��0�Ն�j�<)���j^hq�ӋG*Y$4�"q�<�6f�U��8���'(�.D��q�<��P=k��ـK�(hh��mn�<�%�/C~���m�O�����kS�<�RJ?��s��N lnTT��W�<��g��2YPI�K��s� �w�<9���:aǐ�tc�>L��Xt.XZ�<� ���P�����6.�d���"Om��9s���"S/Tt!�F"O�`	��^�55(�����~���"O�-Ո�w!8ᐖ/N h&�M��"Oܩz@��3P�\��A�^�B�cP�'2�'���'R�'��'��'
���T�[�qw��B�ִ���'Z��'�r�'}��'a��'�'Txi�s��3��]���C�/����'���'z��'y��'���'�B�'l�j�(�J
�hkR�F�v3��'�r�'��'j��'\r�'�r�'̺�+îW��
��2KN�/�<��Q�'��'�r�''b�'���'�B�'T�4�#K�n�ҩ�3n��=�%k��'�"�'�b�'��'c��'�b�'mj�Т�~y�A��CT�9�i� �'�B�'���'�r�'���'���'� ����+:��:��N&5^�
��'+"�'���'���' R�'\�'!rO6*¥ ���"8L	H�'���'����d�'{�''2�'�(�S���>�"�$�R65���S�'�r�'���'��'��'���'�� ���Yj�`�T�� Xї�'fB�'�R�'�2�'o�'�2�'hL�A��U6��P�H�d,�-
�'���'���'�"�'�b�'&��'��@X���^�����)�('��(��'R��'��'�r�'R۽G���'���H��D���]#2��BO�$���Oh�i�ܨ'�|����<��H�
��R��),�R8�P-4r��G�D��5��7i>b>��ޟ4���3 }́*��;^�-S5�O�l�+��K�3�Ĳh[��䦁2״��Ȉ���>QȐ�VZZ��5�?1t���E�矄͓g��V�O|����ӽ��)\�]=~Xò��Z���s �#u����-71O���d���]5��T!��Iy�Э���>��Iş����*�?�v�W>��'rSN��Xw8�'2L>(�GÁ#?B���gJ�/��d�x��9��+��t�Oh�Ƀ*���'�Re�$b�L��jā����y"^�&�L��.46�lc�(��
��l
禁,��h�F�����a'?�\��������a+R��?9�
�r�f�1��Jn��1����k[��u��4h"�9�rM˸|b5�O ��p��-����iL97��1L�ʜڀ�/&�<��?Q�ltGJ��|���䖏1�b���H\�%���� X�g��$P��1Ox�l���4;�?��-��N������j�`p#�:q�	4]w�Ez"Ɓ�S�O�5o�k��Ώ�4�z�	��M1VO�$ba �$t��P�n"}2��O��;���Of�D�Oz��䟨�ʤK�~�,��a�'&�����G_�r�-���;3���?���?��3{��Χ�?��o��WM���PF�e;
1����.��I&�M[b�ir,�'�z$�S��~�dL�IG-cb����)�mnp�ـG꒳'v7��8%�ǭ8�Pם/!S�	�nn��
�'����H
�!�\��G��K�t����:�b�'J��'�[��a�¥Ӹd���3ʮd#��3���� �,:j�=���Mc�[#��'�H��?�۴Fdj�[�*BSr��b�ЎZ��a��W�C0l��2��<��rc�4��
c�M����Qy����s��5SfQ���>��A�2��[��?9��?i��	�\��O~λatlt��'݉,("xK�Af$9.O��$<�҅��?I��4�?�5�j��	w0a8BǄ�F��HPsN�W�ꕘe�OX�S�C��)�V6=����z�5�'�|����.u�v��B��E�ҩ����:����	!fl`�jUD(���}��:c�����O����r�2��NTf^i;v�9���O��WR���?�?���?���<��(��)�8���\
M��H�a�i~���>��i07-
�k��V��j!۔�O% M�sI�)q.����'RW,���%Ц?۶����
�ʓHS ��'��Of�G�!�>�Q�nC>Hy�&K�X�2"˩-��a��'L�O��'{�3^�|�PC,'��)ˑ�@����`�����lZٴ�?�c�[~��<�شfAZE��^�m)�{g��/T��$�i�R	b��.pک)�'��OU� �T(��vo��J�O�`���-ŀ]Q��ؿi���k���Հ��'R�9�Q�'v��'�R�O�͉�V>QC%Z%,Ȩ�`p�͔r��6�V9K��Qc�h�˟P�I��L�s���'s�7=��⑋I����ő�9��qkY[-���eӚ�g�O��8�MS���ɜ�d����� �D���Vޑ��Bz��Q�0Vj?Iqbc��p$���'�P� �'����'���(+ L�Q'ϓ#����=k���'S��'o�	L��K�Ο��	�q�N���8����4��'�۟�QI$?ys[����Ŧ�袟����_�I� x��j�/��15� $��D�O�̺��{�hrJ�y�˽q�����:��ؿE��D(PA�0���A�T(�?q��?����J~����?!����J�Ω,�:�plω)'�$��:���Γ��DW����	=9��Ӽ��KgǳK.����&��$1`\�
�iv0�@G�H��|�\�I�l�*�������G`)��΃p<���0�\7O�l|�q^���q�Ɵ�bh]͟��	����?50��5t�r`��H5F�da�ĩ�<͗'�4�Y�V�p��Iş|�s��'��!BFH(4�~��E��
 *�\�\�����vM��DIPm���)쟴U{��#Nn��'/��(��ٺIO1�p�Iy"n�j�4�/��iϸmO���Ь��Ju��anH���j`�3�5���$�O��d�O���<A&&f�����gF"��*��dj�pp!%(P��h��*����'��O���'��7�צ);
�=�p�v��"R�F�;���$'읺��	���x���g���J�����M!
�K�~�����  �f˗�g�.PPCi%X��5a޿�~�d�O�D�O8�i�[����G�"�.tE�it�Tnރc~���O|�@����16�*�$���-�	���ɕ7ANh���eֺ�r4.��_	�My����ȁ/��4��u�dvݽ�'U\D8���cz`tGe�Xh@ �.j%�	|v �'�^�D���u���?����?i+Аw��9����09��A��?������@�x�̉)�+�O��d�Ov�9O�acr+T�Z��D	3��C�4Xǜ��;�O����OJES�O�d�%�	���N�:AU��ɷ� ����Lk�p���J'u��(ڱn�>�S�V0��?u�A�`�
Q�M�6`\�QE"5bv�'w�1P*�2����'��Q���3�'B�Ĵ��!�\: !Ǎ�7U���������3�M{�J��'D���?���7=�-��i��MB���^��?	�N�E ��sn��<��>�����dݝ�烀\}r�C1M���!��C��L�#��?���'�����'d�'b�O��mcuR>�z�$�šw���QyVQ�f��X���@�mA]y��'�����t�'ʸ6=�D�͖+K9JQ����j{�蚱���y�4S�=��3)���!?ʐ��u�=OX��6�Å5,�&P?[�ЈQ9O2Lx�,��y��r���ßT�"�܉�*����tȣ��Ֆ�|9#,J2T����I��	ß\�'�T�2$���'oB�L%>�$��i�9G���kƯy��N���FI}�d{�~�m�z���I18�P��O��<�gŭ$�}2a����Y�t�mZ7a��'@!f��r��d'�c�m@� G�e�s�C�'#��']BnSUj������'?�'��ŚDE]J-�8x���A4ްZw�'m��Þ'�R�'�7��OTM#����]* 0� !���:�|��JQb���ڧ�ÃdAⰢ۴zU�����Ƞ�u;O��!w��]�M��T<X]L�QA� �:-D��/bx�'����;V���$�O�D�O���ũ9~�Zb�
�lI�#�� 
t��ԋ�<9�F�7R����?1�����|2��u���+rAD�[cx�g�m�\�3[�\�4'��Mܬ�~�k[?j*a�����%���t��䚌3'\1��^�B޴Ih�!r�p��me��	��>�'���$=D�|%�A���Dɇ�P�8w6����'^r�'2"�'�剝=nl�c��<9��@,-��ZDdE�4�(�ـ����s�4�?y���}~B�>y�i�46��1gM ��@��3����O�/u����C�>o�j�V8OX��X�$=2��Xw��:eW��;a�g�н(�8"��G�4)̄J��;R|4���'U��'���O#�Y�����w8���/ƨlϾ��3�Q�I),�`��'�2�' f�#�'8�	��M��ah�����)Ä��L�I��E�>�ـ�G�{?���D��uK��|�5
L���'��s�3j�u���N	��ŋ60��I�r�� �'�d�$��u�͕��?���?�¶(Ǡ	Ee��>���۷A����4�?9,O����LϫA���$�O��D��
7͈�+�2X e�]��<}�@E�2xL�/9��
�M�W�iD��'o^����|*`@N+��Mc$������`R* ڌ�AC3GSr{�S��IФ��J����I�5�4X�"�pU��#GS?,�d�Z�	�Z�P(�&�?���|����?!+O�0�@�^$sL���l�$P\d�&IǱp��d�<I��i1�	ʹ��DDf}�Gm�A�շZ4Rq�v�H�5�13b�Ԧ��6��@��ѥ4?)��Z3XX���.w����'����$�VX�hq��Q?9���X��L�&M.����'���'y��e2q���$`��݂`ڹ"��Ef�D��b
#�B��	�����?1I�yy�O{��.�2Ɯ?"�pg�6����Mu��o��	����=#�A�S�?�W�B(mm�8��-
�XB.�Kk�At���B�ɍMP���'��, N�����c �|Q���?a�j�"��7�D0~���W��?���?)���d M��;s"�O����Ob�����36��8� �e�˟�~�2��.��dz}2�a��=lZMP�	�=�2 +D"ƴ}}�Ͳ���(eҰ���'o�/� �����xS�L(�R>�����O�9AC
Y��ipFͳ��Y�J��u�
�p���?��9������G0��'�?Y��?1�Ə�FPhh��GD9\p����?���C᐀a���?i��i�؍��4�6��aՇ.�h��#�$>��hS&�
1��Ϧ݊�k">u�%�=?��K�ם�k����эMI�t�AIέt��kq�Rn�dMܟL���埼��П��	�?1
�I��U���aRH�;���i�T�]0���'��J��'AI�	ܟ��s��˟�%E� �d@�ЉS��A&����V�(�40ɶ��JT{3���?���v��BЏ��A@n}Kb��
��� ����J���"{���f ��k��V���ɡ�?At�2��°��&�15n�=��-��*��?����?A��?	(OukÂ�X��dގ,(�!7"�2>�5�B�!���$�Ԧ��	��L�)D�	��M�g�i�t�ʥJ!�=��^1t�|PIP7P�� ��i�#�yR�'�>U E+WٺS����Dx�}I�;S�n*u�K�XL4X!���x���Jw��M���'8��'����{���y�^��20��Öΐt� \[���'C�ώ�?1�O�RLa���$�#��D�/�H�HЋ�r�0|	���5PP�����O��2��pɪ7��ఢF�P�r�����O�e�oQ�[\x0K�G�:ؚܓӆn�"���vb6Y�ONT�ɪ�hn�:�?���?��oW/Lpp%�h���BU��?Y����$���`
�O���OR�9OZ9C�el�|��Đ�	��A���K�OF�mZ#�M���M?)
N���S�GƁ;R��Zhc��P+)<£A�TU�P�
�S2��8̋��'���CĲ<gELi����D!j:���h
�vB�[F*@��&�'��O,��'O��~� -x`'Ƴ^"��S�W�q��Qap��0��ܟȪ�4�?��J~�c�>鷱i�f�; "#]#,l�UnH�.���T@v�"A�E�8�ܭ�U0Od�Ą,] H�\w�tmіY�� h��E+�&Qt�!X�{�Z�:�'K:����U����O&���O���]	c��'L@��@�܊;-��7�2c�L�H�Gד�d�����?Q���Γ�����]��^524�ݚJ��$
g	
6;��$�ٴ����R��~BLG"T�ON��!B��,G;� ��[���
p ؠ#��Y�Ep)ΓD�J�AL�O�� �>@�'0}�r�'`�B�!��I�`ܘa`E�󆘺*��')�'J�I.t����ÀП$��������ʷ.XZ����%HR� �!��L�ծ/?q%U���I�Q�4��Ȓw	�p�p����=<$p�)�(����<rpR��^�XsK?��G��O��df�8�ڹ*�j�Y�6�����`�����?���La@�hW�Ў��'�?���?���-����S!����3��֔�?� �G�<����?��i�Jӧ��4�#��J��d�B��;���p��Q���`�-�����_#3�	
F.���I�Ph���q�'��fP�)h���'��Qs떣;[��'�,��I���擖RA� ���զFK�pJ�h֮��Ih2�1?iu��	^`���?����S���	&|����0	=J%�����3��aJ�VJh�z0k�OV����_���iQ�B�2����A�{ad�:hˁ8�b� ӂψ>���']���Eڟ�Y3L̳��ğ� ����mp��kV1<Y� ��N�5!�,X��$�ԟ��	ڟ���ݟ�'Y��� ;"ub�ɄtB�X֣ņ$��i�(H �y2�v�b�Đ�n��	�����)�4L���̙�Y��3U���#nY��fQ="?�Te�KU~ҽ	��4#^w�S��~R �wj����G�X��Xsq��:�~�`wH�@}��'Zr�'G��E۱.���ywOG
��d��喎Y�a�C�^.���'W��X��yr_�@�4�?��OV�<	��X?V�z�-�� �`�h���$~���E���;т��M��'(��ҽ<��Nӟ�$'���ģ��s(��R�Dh�p���'���:H�{�b�.�]��$�$�O� 4i�\���؉7�.0��zcX�D�O�˓N�bP�AEƁ�?Q���?Y��<�aO�V�t�(R��f�;��W~�l�>9պi��7�Էt���3�����OE�DbR������˙N�XY��AM	&z�,���]���	���u7+L��?	dF�d��	'MB�y mʗ~h�`[���$��	4��I稇��,�i>���ן�'�H��C�Zm ��+5�A?PFmI4�T���	�6P�\�ݴ�? k�u~�e�<�ݴ/��]���!4*Y���D�mq� �i2��Mį@�<�ĭ#_¤��i[`|��[j�h��O���W���\��4�U�14l^y�`�'�����9F����ӻ}����>��f&*Vnt��V<(���91�� �P����?������Ir��-q��U�o
>(a�+�.��IB�K�`lگ�M����o?!�_�v9�'K,�	K��ӟ$Pׁ�6��}Y���"U��J��O�<�Q(Z����$Ot�/(2KR%�I�q����[Y} �S��J1~���΁4�AQ��O����O����N�8nH��f�9�(���OVQz%��@�O�TnZ��M#�ǎf?����0ɘi�I	5Kꜫ��G9""�h����KL�sN�9Ԟ~R4�ڟ���O�DPe���Q|�(�&��-;BX���'��';.8a���+��O���'��H�O 2UXqM�U�N�	�hL�2�"�T��y��'��q�b�D�@b����Ɗ��VF�L���W�m��I���mXf�Xsm�=��I�y������y��'�2�� +�5���9b��]��K݄e$8PsI�xצ�rL�����V���r���?����?Q�'uĨU	��X��PCPn3�b�#�M���$�6Yl����<�����|"�[_����G��L�,�r��M��S�T���ش՛��I��~Ҁ��_Y�H�O�6���]�f�s�)�Hg�x1-%n.j�5�>3�4g:��O53��bd�
XO~�,N4ld9�#�7�<�����'� Ʉ�ɗt�]����ҟ�k�a�$R}�U(`�G�(�>d��Z��T��4�?q���m~≴>q��i�87mweh���ms�ASh\9���B���$�$-s"����  ��V��N�[��O�l�Ν	\,����@t_%P�� z%������O����O��Iޘ�|���F,��3�LZ�F$&AcpFY>sn���O��ĕ;z�<��i���[��y���Uw�h�Jۆd�I�$���bYs�'���k['����O�p�[xlHߴo}��䁡c�H,vkȻ{׺����Á�T��$�Ǔ�?������WϟȊ#��p��'���' ^�:�l��o�r	rG�̾f�����'��X�(KS��ID����⟠�	�?7mHP�� ���_�,) �`sN�#)��P�'�~�9��h|��%� �O���g��r���F���@t���G�gZb݉��z4`Y��D&V|$Rf��\?�Yw褘���N=�J�O.���R�:"7i@��@��K���a�Ε�X�v���ߟ�՟��Cy�hP&�B�2���%rh�Kti��~L��'L�6��O(R���êO(n�4:�m��|}*d*����⠱�4@#�M��A�|Xoڶ8Sb���i^�ݭ;~* D*��O*d�d�s���i��25LƜ($�'���$�V-��d�Op�$�O��)�i���'A�XVc�)Ue�t�S��=����%�<.�h�I��?���nھ?��	��Mϻ>�8����h���m�+| ��W�i�p7m�������c�p��F�Oy�D��/J�@�ܴߎ�X%�^�Q�@%�_�#�����5O�U�Ю��?��&Ϯ��Dݟ�x���v��'M��0�`�7��̓��E('8�e �'E��'�RR��i�M  uф�']�)��Na����A�D�b�\�c�����]|}��'|"
���~�#1@��1�#��B&�)<�L�+��W�j��	53��
I��^���h�X�;�@P�I�@w��t6�3t�J Z�69��#�:���'�b
� ht�58�����':R�'׈P2�OL,o���i@Ƈa/yZ��'��,Bjm�����O�Hm��	�e!?�;I� )ۖ׵}���s*Jj���aɎo���>�&�!�-F� ��+��<�3k�� K`�](E:� ( ��	Ҩ*�,8�C�8y�V��� h>剱�?�f��M���'��'���X&K�f4�J�$����͒�a��$��Y�j�l��ﬕ��矴�I�?���|���l���D��:X�ģ%▮D�pE�B_���	͟4��A����s��4D"������[�T�e����h�0����Pj�0'�~A��O�4?�ئ%Z�[�����CU��:��FqD�`l�jW�����H�q��h��NY.'ӆ�*���?i���?����:|xT��G�O�0�m�:kg詫R��:/ ���bj�O(�o����{r�0?��^�$�I̟�a6/R�%=j�Ig�� H� r���cB1���% �����@�$T %8�Ƌ#�f	��'�������1� ���M�,	@��ցRkީ��i� ���O���ퟜ@��*�9�b����
<i3�q ��4"XWo�<i��hU���T�'J6��O�x�6O��{ץ�'x\�Qf��/l��p�<A��d�)-8b�'��iݨ��(��$<S�b�ȯ.�6AS��5|���M���B�NS��ts�aݫ��������g�ǦuY��?q��:�I2�
[+k��ɛ��|Ai���?Y.O.�7o�)i�F�D�O���䟞Ȓ����cn�5H��X�Ew�|w☰9��I�����ucش{���7��U0bim>��r�-��mjER,f�D��B>@@53C��?6T�0�n����2=L�� �P��H���]�9�B��1<g:9�Pm�矀s��(h�� ��ٟ�S����Yy2	T�m ŏq6�111é�0�K�p�H���O��mZ�� T*?�2V��	ܴ/o�s\#V��hW�cC���a�mӚA[�鉴v�1Y��0f���Q�q�d��_wMܤ����<�dF��+��̱@�ԁ6�X6�K̟4���[�lt`��?����?���9�z�:/���;á�"Y��(�B~d�jq�]6Q�xU3l�O(���O������S��j�����^]�ѹF��~�|�a�L^�?���i4����c���[�%#
��D��m�.,Mb(C��w����ÁS�h�0	ʤ+a'�O(�1U��{yZ0�d�ON7���<A&MZS@��	'u�q(�ҟ���ڟ��I\yrDѪ8%TuC�'wr�'ʈ��Ă�3�xY�L��:�hѩ6�'ƨ�K�O���'F��'��u �'
�l�^EpLh*`�,�ri�U@E�@�:����O��I )PYF�[��غ��u׆��?	T����49�B$���r4��)N��35��O����O���S�+wٌ������O��U*�D@Q�R!F�`XB�-�H�䂛F�.1n�̟��Ɉ�M��R.���yG�Y�I|�LZg*ŝ.��U�a����"s��A�l��$�Y�0a�U��'@԰%Yߺk�Ǡ@��D��2�ҕ ܔITZ	j�<1��'V��30�i�x�D�O �d�\��	�6�(��B�T�v���>t�˓�l��"@
6X�-���?A�/�IB�p�L�<�jY�򬅍\f��S�傎�M��kP�fw��-�SL_4Ep+S��-��i���� �`ß~Le!PC��(���n�=x��wLS~�@}L��� ��~��25R��+��As���BO�u�i��QCx�H$`��oy�`��?��?����$��T���
���O(�04�-HR(�V	�m����3O:�d�Oh���5O,�D�<�ƾi ~�ɇ�{����<95R}�F= N��cAK��\.���U�C�`��(�e ۋ?/X}��'�n��}�DN�
h��h�gMP|蒦F�am-�?���?���:���bK~��8����ޫp�h���Hެ1A�Ap���?a��p� 5 ��i
�������)q���	0+o.4��M�Gǔ\���4@�	�b�p��qa�7%���4�b����V����dM��?!��ԅZEj@�6��kܼ��`9!讙@e��O� ��Mhy�m�O�C��O��$�Ox��ŚI=� 9}Oy��F�We(� ��'u�l(�P�PQ�b\$'JD�Sß����?I:ڴ!ߨ�zg�'p�BX�VkÂ����?)�O��{���j��O���c
BYa�� 
WrГ�'��#�DK�厨WJt�sU��1AV�\�p&���y����L�<j���/�<qU(7	���Z��j&8e)�6&�r�ʀ}�yI�'��O���'E�	�+��pA��]��� H�S�4�fP���!xЅ�I��I՟<٤�z�,�	my�Hs��;�l�0|�l�㨘�hMT�ࢎ�Vn�2j�A��J��j����Ig-&`�"�юK���Pƥ|�����15�N�@E�Q�k�z����O��4T��ش^,��'�r�OQ&�W>颒�����Jb�P.��4�&b���fNBD�b���O��d��& mZmyby��nޥzw:�y �C����G�E4�&XnZ?�M��Y?�fG�)�����?(�ʉ .hl)�'Z�v�~(�sk�=zH4����'XgJ�M(�K0�'_tX�vF�<Y��'F��q�iR��ĝ������	���b"�-�����O��D�O�ʓW����1	ֱ�?!���?��K#�8����xPih���,�?Ab��C~b«>A �ix7 ��D/,� � ��;��X򂗛d�5��fW/�yRm�%9�x�5��e��)�h��#�'�RI��%T�	0��a!��t**S�Y�	ߟ����M0D�*�F�꟠����8�' OD�ƈ�f�F��V������
4�M���?)��i��Ӏ��4�ؓ��	W%NA�S��)�e��@':l���զ��Si��X��'-C�h׋�O��j$�Y��ugoنCԈ�p��	^P8� G�yj:�2��iy#�Ov�0�x����Iß(�I�?Q�����J���I����1{$Nǥ�8��'cD,�d�6X�r�'a��O@�7=�����>4ƚbP�I�,��$CڅMe���'>6�Vʦi��f�����C�U8�����*T��A%2h�WL!"�܃EH�n��t؟s��I.D���@��A��9U�@���CI)G��;V�5��ǅJ�!j-���^�?1��?����?�-OV�Y��۞7���d�h+#�-Gg�l#�M��;�B�$ ��m�I!L�E��I��MS׹i)�HJ��8��Q�m�18��H燙|ȴ+�. �e� �a�':@��e�Ϻ��
*N�,�IϺK��w�Z���t0���e"�8o�u@RaR	O��(�Oj���OX�Ɋ�-F���� H�\0���LK��5}�&���O��ėX�JAoz>��	�M���-�LQ�~
|���NJ��}h�N�..���@}?YGk0D���۴����e�ε���?����y�? �qwAI:f64�b��3!�~��Teu�ك�
�)?�*�?ɳG��M���'���'��D��ҙ!� �g��y�H����'��`��Q�����l�$��ǟ��I�?���4U�jlQ��l�Y�K�z�ϓ�?�.Ob�D�O�� �>OJ��p�Y�D��;R�>�I#�>.�����j G�(��ʋ�7G�䳲 �6\�k�AY2Mm���KT�p��'��� �c�(^���)��\��x�Q��O
M��g��0��$��n�TY�t��O���O���ͅ7$M��P=@������dB:7d�u}��'i"�'���'�(��d�w&��'��@{�A������w��c��'^�H�1��a�v�I�_��a�+���b�� X8�s�'_Ƽz�5�@*B��W�p�H�	�����"�?-�Mk���P Q��i��o-����_^$jQaV@�X��#�h�$�����O��d���Ilz>��I�Mϻ���吷n��*pJ'A�F��W�i�6͛$f��d�C���h˟���[�QH���We��[դ��'U�/w����M�r���A�bAٚ'oBl�Z����{��8ٴ tb���7��0Ņ�<7x���2gт@���'���'N�Iz���ՇU[yr�'ev��4U,#l0����;%���[`�'�H��'��R���	��5���p{P̊~�ԙ���D=��z`F 4a,<�ƌ�O�0��#�f5nDCƄC~��dh�	C��O����;A؜Á.Q�E���( ��+q��\*���?a���z	*�ą���'�?��?I&FέW"Ց�i��!e���E�۴�?9�Ə+;���'�"�n�L���`)�iޡ1�k��y3��y�Y�|� �fO�\hh���l��MK�ђA���p�WrL��WA )�VM� �C�U�F8�D�>y��׏~��0Y�Y�D���}�d���4|b�'�r�O}�0c�IԼN�l�[$",y�����L�`��Ʉ{rV�������������M.O:���N���	 !(�;(<���\}�
`�r�o��p�I�vJz,���?� ��X�8Ş4P�D.b��l��{[�U����e�4�I�7�ҁ�'�'�z�pJ�<�@�'��8�B�Zl�^�q#ד{-��!��_�^���f�'���' B�'��	�3m�@R���韴��N�CZBQ��m,����l�۟(��4�?a% A~�>a0�i�6��4'���P&��:�h��ԭ�3@�Rȗ��08&L ����Gf��U�xH���XwI2�sc�St�dK��~`Ҥo�8t�:y�R
Y�7��8C��"m��6-���ҟd�S�.Т�&?��
H��9h$%��u�n��6䕵M}>��IßX�	�pe�U���|z��(��V�'|�l��'2� �� W�D�#>3����A�"�~��CD����/�Q�F�w,���y�!Î0j�I���:�<��F���I^h��D�Ɵ�y�ů��DҟhP����������?	��hy�-�
������p��?�)OX���ܶ�R�$�O(����Io�[Xmg�љj�ƌ;��̮E0��v��Ɏ�M�Q�i�ƙ3�'���1�EF�|�)��h��Ye��8G$�L;>R���	3P���1	
�<�S-�d�9>�L�'�Xz�ʟ�L������>1�tD�OvE��	+/�����O�i�O��$�<���՞;j�ࣣ��V��[�J�0j�%�Ӱi��'�z7��O�=p��Y-O6�O�;�6���ƽNҺ�bF'w���oZ4�����,؆�I��~�|�tk��y����58Jȹ;�')l�ň��X릥 ��� R���%��aQ!%�+�O���O�����T�'�ze(S�{q��0��˫N8��`�'��H���?����J!�����'�\6=�j$B#ㇲh�d�@C��S�H�j���� o����	�lo��������\5���j�-��_�dE��� ;.y��PDW;y���08O \�r(Z��?��29�	�?�A��M�@�'�������*}�A�>��XK��'^"�'R�]��Itb��\�"D������I;���QIѵKߐ���怓c��i��Q���b����M�5�i(�u��'l��Q�Z�*=��0�*�8Pd$�6���0�:Γ 13�m�_2J􀠌�Z���O��?�-���̚�f�*Ȃaȡ�/2��܈�N�Oh���Oh�Qj?dﶒ�6���O�.H�\������)�b��U)I.@��D7�plZ͟�I��M���I�:��)�����u�僯|����a�L�����KJ�A��n�#TřQ-�7�H��`�٦M����xqk�'���Xz���H�u!O%#{��MH"�������OL���Of�	Z+
�����e�y{�ILl�R��<1n֧_5ؐ-O�����v�lz>���j2.�z�̈5��˕ʢ9�"��O��m1�MC$'A|?��I42��ZtL�ɒ9?N��%�͛@�x i#�"�,!uC��<!���/9�0�	u���'@���\�M*��m�6_ŴI�`жP�&
�� ���O����O*��<�Wn@�L�|��� �t��B�N0�@A��:,ll��t����'����|�t]� �I˦U -�T7d� s��<@�
�[�l̜L��U�r朓7���D��`�D^T3��M<\� s�'#��߹�B�ʁTa;��Ȓ���D٫f+8lڛ�?q���?����\�aN~λc��#�	_� 4)��:�6< ��?����v��#���$�'5�7��OX�1r<O�HX'�Z�{�Ԥs��V+�r�lI	��dJ�_"5&u��K�*�V�s5�B���	�qcN�!Ƃi�H0�H
Yj����?�(׆�-�?���Mk��' ��'9�[��]�^�n�P��R޸-��'EB\����T5~�����$�	�?E�ߴ!Ⱙ��0#��	�i�,��'�x�"���fdӮx���O��+��B���t��'sRT 0�x�Z��E�޾Za��s�ƈa����]��y�'X�f���&4�-O��`�/A�)���@�>��b
ğ(�bDI�q�Ρ��ޟ������Oy�@�9qa��&\�I���ۆ�:�aR�~�����O��nZßp	0�(?�[���4q`½sdǖs��X�T�ϙ0|�&�i�
Ir�O��f� �"�͓�y�h��w�᭻ ��$�wO`�D9�ō����q��W�&�@S0o�O"�I����o��?)��?i�'`��9 .��yZr@Q�����)>�zTA3(&S�S���O�$�O��I���S����ke��3?�Ð��%O3RAu&����o�4�!��OHU�wI�����'%�ʙ���ZB�� v�[p�܂t���Р���"�����7O���A���?Q���ol�I8�?��2�Mc��'���G⛲k�m#�O�UkD(x��'��'��W����lm�l�	ߟT�IJ��h�쓨[�씫&ǅD|n��	8G^F�F��	(�MW�i����'���BCÉ��v�΋ʪ�0T�\���36��CCC�a���c�ȉ^�TL
��?1�(��p]PDFC�U��9�s��B�I�v��O�D�Ov�#��U�@yJ��L�D�O|�D̀-Ld���"X>�1!�%7���É�n�����I��M���*�H�yg�]�#*��Dh��c)� Z�
K;6(Yo�Ca�7��fz���e N�*�b�jT��OH�£'��u�.ȩuĬ��<���$o�5A6�S7�ZJy���O P�%b}���ϟ@���?�"��0��0Pf��N%n	Ѡ�^�3��-�'&D��EB:��I��x�S��M�'�?��dM8t1�&"��<���7�	ڟ�nZ-hT��I�$�,��q�?�Qf���g����$5����"�(��q��/3���e����2OD̸5�<ɗ�'蕫U����+#��q��8��唞nH����'��'hR�'��	("�J��Q��ɟt3I>L�����/�`7
���q�4�?���E~B�>���?�f�ĩEp�Y��J^�)XimJ��)��ͫ �<�&�D�	Dz�]�BI�� �P>�2��m=�� E��O��sb��Xxjx3S�I��MF�'y��'�����g���yWBS1S�b��V��|h*��$� 'R�'��e=HMP7=�h����e��5�l���� qJ�) ��u�R5
�a�F���@�Ȉ<A��4���#��G�� ``v?O�4Y�ۭH||�ff�j���
��V)�٢��d�P�p@��"��Y�4 �b�'�R�=�c�C�v��}�%U����'�	�K�f02�ן0���X���MK��^6e���@4Z������<	�62�	'�MK��i�$� �'���8s��|�6�P�I@�Y�Ϙ+���"<n6�����S�D�<�� [R���#�T��'����eƝ}ʰ4���+@�$��O"�Z慂C�"���O�)�O��ĥ<Q���Q�PH��d^��G�ZZ!�=U�iR�'e�7��O"p�Ր��#�Ob��ـI����NEkc��8�,�$i���Ѝ^�� GaG�_����8O�j���u��V1!�P̓g�ԭ��-��c�6EYp��xm���	�?9D"� �M���'���'����7��i�H̋�"��9�HCv���8�`���S�������I�?���t���l��N;�0��(W;��`n�)F��o��Ms�L?��Q�G6��'b���e�єH��SE�6.R����aJ�,�)���<�r)� V��4v0ė'}T�d��{a�7-�ϟ���,�����FH9.Ƶ1��@ן��	韼��]y��Ic��b��'wB�'�@Q��U:
���$O8�Ҝ��n�O*��0����-O���`��@@��O����jK�7�"<4HZNQ�����pØ'�.�� �X���hg�]���i̅X���������V�ᡧ"\�> x��nT͟l��̟�@��A%֠�%?��������$W�U���Q	Dx��6W�^h��qrpA�4���I�.���Ӽ3���*UX(Q�EB�T�<����� �>%X��� ����
�fE���'����Hߺ��Ӟ�26n��#�e����2����I)��D�۟������A ��?a����lIzɘ�X���5\�-'	�U3�,X/O�(���R˓�?���L��O�bB�,L`9����&&��9#������f�jӠ��v�OF88B�{�T�O5H���0IJ0p1+O4m�C�"�?mb5S䢞��y�f8[����00c�(�,O�4���w���Ҏ�<)�p�32ၝ�"�ᘼ�J%�����⟼�	{y�%�����'\�8Rb��M�)vᵬ��]b�fӎ���Fh�I�����O��$K��hU�G�y��(A�+>��ҡA� ��flԷzy���@Q�_w��+5���<�^w j��K�����TT����+���jd�y�|@�	ҟ����?e�e��Y�sީم�b��{���{E*�#ڟ������J�K��M�Op27��O�![8O��3̋�S�>E��g?����''M1���[%E��MP�����lI�eΠ�KT���y��a⺉��4~8�d�ǊF
FL�1%���hÔCH6��$���؃��Φa����?!���4�1��4S�|9��I�u���?a,OF����A�I�.�$�O��D�poZ�����َb���a�me��X��I���l� �j�ɵ!�n�7;��űQ�V�A�nlP􇊚X��&����J`���B�ڹ �8O����-�?Q�8 A�I5_ �a$ϴ\V�=vI���x�	��\C��J$�?���|����?�,Oy@@h�6M���a�W6�$x�-Tn4}o_yR�b�N���* �������T�Q2�!ɐ~d@g�O�GHQ�-�M"���p���H��͓#�\����m	6(� <�><���;$OݾN����b�����O.�{v�n�,��I��|���?��S	B�T� d6R�+A�&鬔�2� �f4VQ�7�8|'��'O��O��7��<A��y�O�F��AƘ���a�ũ]@�6͘�M�ͪ�"G�W�f�������A�SI�]��		V�z��N�j�g�!1����S��@��!�|Y����s���ٴX"�L'M�����%�:;�p��c�[9��'t�'��&e��Ȼe$���4�I͟�p�C6B��(b��?�� G�SʟX��,?e_�|��˦��s䧟�#7��0�<�����c�H��������P��/o���C*`B˧H$����#�7�V=&�b��C�,�h��4�ǀ�"�'*�H=Rudta��T�'3"�'A�Up +ț$�x�x�U�5��L2��'��d㡯v��D�O��o����Q�)?ͻ��}���Z	4� ��%	&���fV�3�@��i����"ZHK&�k�Q��y���,R�;I��ɘ�N�ń�aW�kP7M`� R\��k���40���'d"�O<�I�▴d��cAdK��0�$�Z�I�2�ڤH���џ\����
�M*O2IST+D�d�3�H�5<��4Kq}"�L,m��c���I Y�8��D�?Q�@�=� d�Q��u�DU��#T�1[gg
&b��Y�6OJ����3�?�qƔ�U��Ɂ�?�]@�^��$ C�:�BɈR��!*��9�M��?A��?���?�.ONlÄ�0!���K�R3P�#a���"��T��A��ĕ��9��1'A�����)�MC@�i^(�P`HvD���O�,�8��Fת���q�AT�`K �'�~�فiѺ�gI� �I�#V�w ��PуJ�L�hXЧ�#��hٰ���G<��#�O����Oz�)�$f��󮛡aN5KWL��TVTȤN�G����O�$Ê1�%oz>��I"�M��H}&4��U�t��=�M��YOx�)p��O~?�g(E.m����۴�b!�-6<���w�]
�?A1/A��`�2��d�2 �&̓�6�(����O$��&CGyb��O���� p�:��	ޟ��	�C¤5� �9[�cv���V&6E�	˟̗';&y��⛣(���<���M3��K����׎&Z�:�k���k~2g�>i��i�6���~����oX��F�O_*�`�ou�H)�A���`��U��>F7��b�u2�)�'`�n
z���umL�Ft����Ϫ?Bdz�lG�R� �W�'~��igB�#A�������'�^�Ɂ��6i�x�c�6u��d	r�L	�!�4�?���mW��'f�p��O��'[��ѠQ�� ¥H��+�HH+G`^O7-S�Mfd����=��H�� �OF�K�a�$�u�G��K~`h�:i��Ä1Q��a@rƓ,!N���I��?q�J��M�$�' ��'�����T哽fܶd��Ȥ(�RR%�J�j�g�D,y�,\�	�L�I�?����|���h���wT���Q*ܔB�ąKԯT���
E%�O�7�ظS�$�!���Y��O��䂘�j������4S�
ђ��Ff��0bW��5w�ɱ�'�T��JF=HN����
^�+�� ��;P�L�#$e��'�ȅ�k[:�<�r�U��,���G\�7WpyK�
� �tE؀N�j,5ٰ���:۬X! 	�-׈�@g���]
��'��˖��w���gZ� �hH�)O�#O�jZ���ԍq�K�&�1gM2#]p�h���q��ș�	\�� �9�-�\��G���G���Љ��u�z�k&��Nh�'S�?��)�+�hffQIģ��kւ�G�G<Gz����A�j���K�v�R�J0��l��ᓭqXH��Ċ�Z6 m���ijr�'�Xq��l�Jб��&�j�n��qavӐ�$M3 ��Ā�j��'N��t�'����!˷�Pv�Șb%D�},�Tn��l�IYy��G�s�맰?Y��R�l�">t�=JtS(L4 H�q�����y�it�e��̟��b��_������RCe�$0&�	�t�W:b��vR�XYuX�M[���?Y��
tZ������l&}�6 �X�dQ2��Ru�%��ן �&H9�s�%&��󧏝%8�X��u*��v�j��m�H��Ү�O��d�O>�D���?�����e�)2��Fp�e)�Ey�`�F�i�\���'��'&�������'�`g���Ԁ�S MZ���v�jӌ���O`�� YZ�X�'�Č��'	�&ŝ�M�C�R2+��95�=A�i`E��T�F�m�<)���?)�K�Zxyv�S�[��[bK��׊�أ�i�R�`h剟\��8�	� aG�����ƨL��e��1���z��ā˜q*"Q�|@F�r��˟��I� �';h(�R'���!I&C
d�Ԑ�$�f�$�y�-̓�?�ÝY?�S���I'~ 6��L��;t��Rp$�,)��S�P����	ş��'e8I��ߟ�er��%�|(��O��j-�쉅�i+���'�RO:�~���?���!����'蔙�c�F,�|����D�j�O�$�O$��<qd"����O��9��Y�pw~�h�KV�$� �2KN֦9��X��������O��"T���-w���W�D�GFƗ=���'2RS�|�C����)�O��$�-h5�+WU�ͩ��-Q�-�)�DA�:�r�'8,x0�D�#r�D� d��r&^&@�9ҁN覝�'r$�
hӂ�d�O��$���'&�L؀�۟\(ձፁ�Pj�����+@���'����P��[$%�O������ȠR�ڴ�"M�i�����4�(�a�iB�':��O�J�HB̠�'����4�� ʀ����5[ӷi�d�Ȑ���1u1����
w��<�'%�y��pף�(�\�mן �I۟�A�G����D�����'�p9k�4T�@0���'7X*xp�K�'V
�o��$��������O�$�OB0�D�A���!���&�|�b�ˀ����	�Ni`)(O�*�O�r�,���D�.��B� :�jh��,�8���'�l�	Qy2�'^��'E剁|w6���gH �X9�À	H!�����ė�x`��'_��͟��Ӻ#�N�3��us�i��+���c��Φ1��qy�'�R�'��ɉNL0qؙO\V:F�?40mh�'tSnE�@;�$��֟<����ʧ���OV�F�+Ny� �E�n�[�h�	|�&ON�D�<���\V�+����+a����P�?+� ��Fm�l��<%�����O�˧@?]&�\��ѳu�0�2�U�Q;~ a6�~�t�D�<�����Lz/�����O����t�苲\�v���������	PT?�ˈ̓�u�a��O�N��"q����N�<���y�R��9����M_?U���?��(OR��0�	f����[�B(&h+\�:$Z�4ӳĖ��X�)�S��4c��T��o%Ch�`)�n�p��l�kU���4�?��?���t��	>c���N�
����
ƶ6�deZQʜ4i�|l��9C*q�I柜'��g~Bo7��H���(:���$iQ�^?d6m�O����O�i����<I����|J�'�h�nږmy�0 ޹>�H)8 �E�n`���$�S�'�?y�'���@�M�"iz�A��Dp��4�?A�ԍ���E��)e��Q�O��o��$����Ί1`�Y�PK�-+7�O.�I5��0�I����	my���?<:��b� �I��
�b�=/�8Gͳ<1���ʟ����,P]�O*�֟� ����E�9d����#%lt�2�iS�,�	ڟP�'���I�Q�	�;gE�Xh��&$�Ȁ �⊊ R�F͂?��0O&(�������W�g�6ꂸ<��ׄi>���N'F�z꓉?��?!/O�ɚu��U���'���*���c���H�`�� `s���Υ����y����O4K3=O$�'�BYF�\�	��X�P�>�"	��4�?a����$@��V!�O���'��4e�\Bt1g���%AҾqJ�P�<��1�?a�8>Խ��?�'�?Q�5�p�s��7\:�i�th�ӳiq剄m��h��4�?���?��'t�I�d��;p�R�-Ċh�V��3��A������I�w�����$��3��O�H֣�%�U�O -� ���4~Oh�R�i���'���O�� �>�͓t��,�vJԠV�ޭ��ӪUH���iq��OT�h�nx�|��x� 83�oI�=(�`�@ֿrI"��3�i2�'�B,G�W���=~1ϓ�?��AΦ�2�
ӷh�$�:���%{�%"��w�V�D�<)GM�<�O[B�'W�
S*v��y�с��k'�yAN�;]d7��O�H��w}����y��'�R{�'�\c��@� �0"�af��bZ�A�O��P�����Ip��ߟT�'��`�óWH����
�2+Č{ׇK�/><�Rޜ@��?i��I�<)�'�?��P��!+��/i'�x�JY�x�J�1j�<����?A��?�����ޠ?ޒ��'.���Hc�׎j���"�ܨ6_�n�)�h�IƟ�[��a����`��!J���	�ę1��d$���к�O���M;���?����?Y-O´Y&.�n�4��5��.��i˥��/'d�%p��O�M���d#��nl#��?Au��<y��|n�f��s�ł�F+$ʹ�["�}�~�$�ON�rP`Ap�P?��	����Zf��G���Z�$�"XZS��m��@Lҟ,�	> :�����(�'���<Ҟ4y�N�() J�RчX�7m�<Ag#�(����'���'y��
�>��F�O��mJN���ű�gY8<
�����?A#�[�<�+O���C&ĉOLL`�oV���9+B+߬,&b��4P4R5K��i���'���O��Y,D�ϓ�(��B���j<�� �c?P��P�i9��'5R\�l��.�ȟ��E����d�9ˀ.���M���?i�4���Z��E%o�D�I�nTF7-	8p�i�K?)�<L�#�W1hśv�'��[���)Z��?q��8p��$/��&jz�	U�kC��ֹi�b� [�>�h���̓�?!�%@�<�����GHN�0���g?C:��sn�a}"�(�yR\����ǟx&?��艵0 ���L~98��FlJi��O<$X�0O���"{���P���OĹ��R�:�q���ţ=q
�:C˅�J'1O~���O��D�<���c��)�<P�@�w���C�� ��G���J�yb�'��p[�'���'�"�ȉ��D�\I(@���ԓ{�8��ȯX��I����	ʟ��'��t�~���\I��!��	j��,���%�$<��i%r�8�y��ުj>B�'�&���}�+�_�����I���,)���ކ�M����?�/O��ۆjWo�t�'"�OC|a� (
�y� �˄���X�T�GGC��y��D�r�'Tћ'��'w���8ٰT�A�h�p���k�7�<13. 	F��'���'1����>�6��,b1�0��*W/:E3䂖#W�T-a��?���<i���U+`͉O��4��W��|J�L�<7��LR޴z���Jºi���'�"�O�^�y��L̓)����O0_��i�'�@�>�*��i�E�'�X�pqĦ-�ϟ8p��X�B�� G֊5��*ר��M���?Q��Dq�<��Z�����w���ɢm	�6-�BȐq���ʕcȴjCD^�T����'�R�'a�h���)�Of���O
!krD&^�,ѻ�g�
j�� ��ۦ-�	�H��M
�O����;O���<V��k��hfh%�/O���웡xH���d����?A���?y������K,�y�-P}����-Fl+�ŝ[}2'��y"�'��E)�'r���'C��أ1�B�Xb%Y�/xD�G����|͠�'P�Iߟ�I�D�'�ȁ��w>��7�YW�*͒ /��E@�Ov�1a4O&����D�4�D�O`{�=O=�GF
���\�(ҡ�h�,`�7m�O��d�O���<��i��<��OW@��t���=4��$aN,}� %;�d�����-��$�Er�'�� #�'��{d�|�����MT�|iUEZ�~��yl�ǟX��Zy"Ā?\�8����|�f��c���;�l(��]@$�k��d$+�"�'zR}��'��'h.�]�:�б�
�bL��u�K�t�7m�<	�ˎ>_���~����B�U�����[
%���y�qQ��@#/�����O*$#��O�O�yp֞��-�7Tî����⮽��ؗ�M�����m�̟���ן��7��R*�y��P�Iy�Ø�%Z���E& �^7�P-X�~��+�$�"�1�����" �y��C7�t
�j�	*ynZ��<�	ןTcM�����jYB�'|j��4\1�t1 ���M�t/X���>�5(Z̓�?)���?��Eu��JA�b"�!{Q̕�mܛ��'�%��#�<�K���d�	�B'��sU� 8�!���jޠ4QDM�r}�׊�yrU�4����Uy���<� �R��[�Q9�]�EC�&��d�<��/�ן�I��(�'�?��hL`x�����R��z �H�g�l�vb��<1-O����O\��<��E$�<t�ׄ>��l����+c�'�>�?���0Uv���?��	ǟx0v����#�8� ���cM#6=K�����d�Oz�d�O�ʓ2�7��!N5S���k�iђ@:����/�&6M�O� 0�Oܥ��'� � A�>� B$;уѱ_�>MJqᒅ0�L!g�i��'(�ɵ0�`<�I|:���у�3��4��E���i��5O'��ho�l�	�T�0!�Y�Ox�کX��`GϾ'x�z�;��[��@�ެ�M+�[?A�I�?-�.O�8��A�57��p�`Β+:u9�9-��'D ���'��'��M+J|�5�K�>��A���5Q�D�R�� �)��`�Mc���?9����V��:c0O�tٗ쐉Ff��+��xp���lŦ= �Y̟t$��7�6�S�dҗ�Q�^ܐ,��ʃ�bI#����M���?����@P�Q��z���O��d�1m���,P�����L�w_�M�H>A�Ƥ�O���'T��Wm��)R��q(D��:]�7-�O�|!�aOay�(@�?q�5|����5�̀Q� 㰅Ҥ?�p(�aC%��D��A�$�$�<!��?����D�5�:hqG�*���	�L��U���@yR��<A�:��<�Oa��'��HQ�TIBʕ�]c��"Uᜡe >�����O��d�O�D�O��{�!�?E�� _�{�m����O��z�c� �A>O����BC��Oz�6O�����M˵m��TƸ�sÔ�!x��sǘ@}2�'�"�'��	��9)O|����a-èo�مh��,ۛ��'��R�=O�()�On=IT�;�	�3�h��EƾQ��}Q5N�@�L7��O����O�� $r�|���O����Ov���  Ox���F	�����2W(�����O$t���'>��n�!��;�Ӻ+�#�&F:2���=Рz�MĦ��	ǟd�1�ӟ,�I{yR�O\�I:*��Ar���@���$b%I�8EZ#ٟ�ΓtCH�ice,�Sⓗl��Q�ƙ.qތ�1D�_��6M�N5o���H���x����d�0����PT�����Ф*[p}bCgCh�L6M\'\ �,�Č-�I⟴�4��
U��M��X�VVd�2���M{��?��������?�����|��	Enڒ;��Y�Sjج�L���Ȗ��b�B��D�s�S����	ߟhEO ����(MU�Y���H,�M��R1V�ڒY���+�O��d��8��s�]ࣂCv�҃������&��t}�%���'j��'a����9�g�2h0J��Z#^%�d,N����4��<5��П$�ɐ�z�'�?A��D�$�(Қx��ꇎ ���j�@��?���?�/O.�� �K�|"5�d��EIˮ�
	9P,�៰{���Ov��R7w���OG��'�nd�O���d�,N��(�߄o����Q�p�I���Ily2�>m��=)�&�h�Ȑs�ܺU�IXՋ�Ʀ����bc<�I
6��$�O�DQ3�d�?*��j���i�Z�2��	���'b�����Eߟ0�Ivy��OnTd����g۴*Q&\�C�.<�#ΐ�~B�C�?ɟ'�뮎�k0��ݣ
�H����K"d��=1��*,�j6��<�v΅0�f��~����rQ�8��@�H!��P@�X
�|�������k�3��'h�dv`�ۜ�{5G�`��@۴ �mP��i���'B�Ox���E�I�`�ݲ�L��yy�L��䂆K&p��4F��mGxBK���'�O�dhT��t���=�9�����^��6-�O�$�O�RpE�Uy���?��4g�o�%/G����Y���ݩ��ǀ]uxb�:��:�	/I����
��<�v"_k��U��~��$�q�<y����R>�	a�$NDv��l���8#�_�ˡ�  X��0�6o�N�x�ʤI��:��aQ.2����%�6 �Z�2��<,	>��C�޶eHj9� /�05�pbQg\4��ju/&^$p���&g4��^�@��B��7YX ȳ�V�T�%��m�,J%t�!��Z�
��"Ҭ� )3�ϑ ���n�Fl�(�BN��?���K���D���?9�O��"�m�y
�#�h��е���GA\��J�"o"�E�E0O���R���@��U�U��p]>��4�Ȗ=`��QL�{M�!��	)#<����O�˓O����;�z`�C$|Na�<�ߓ\��Cd�(��|PƨUQ�.��>���~2��(nc����_*�<`�W-�,,6�ϓ�򄏌9����$6O\��|�u��?)���8J�ΝS�d� h6�u0�k���?��(؉�W(4�f���&�"M��'L/�: l��|
W�׮{��A�	E�]64j�j�dّRҲ�	%B2p��@���#ҧG8-y�@�	�aAFC'���O ��7�'�R�ɟD�h[J� �Q㮞4_x:h1D��P���z�j����� |t�X�'/ғ\���Y�<����6Dr� ㋼T�>����z�V�	ߟ�	����O������0�'+:}j'F�A�@�vǁX���ɲa^�>N��OT|�d�����uH?�OđB�� e>9���gd⡑0���O���������K�"��)W:D�,���O=�� �����'{��OEў�s�þx��4�ժ��uV����%D�`p���1L���87JK�jZ�z �d�.�̓fFx�'�y�[��S7�P?�v��s��6�8���5J��_̟\��Ο �'�z��aC�O��$�3ʴ@�= `0�B�L,~d*PU4����Ɍ�Z�ңJQ�v�Dr&,[&=�$�3����C��q��gh����Q�tM�i��Y �������	8�M�����O��P��""���(��C�W��Y�"1?����W�S�? u��ݵ���T�ɔ�Q�h1�D�Ml�@y���Ms�L�Od�$���h C=s1�<at�>��$�OB6-^������|J�`	7�, �o0?i�\�؊�	U�;����Ov8�,j5aZ82��Xj!����%�.2TE)F��4$�]��n8O�T��'}R�'��GRs��iڀ`�"ul���i�Ux��Ɵ��?E���m)��X�1W�pW&�!��'@"=�ON��P�AD�q�i!Eg�J��0�FB��,BZ� 8��֍{�����O��6�O2%�qn�iQ���F	�~	��z���OF�]{:96�-B����R�	ݟ�I΋U��H#�<�Bb���u*ՐǣR%=��jp�>1ɉ�|<�
���rI�Ż��	J�$d@��i[�/3�D� %+�k\���	��D�d�'Q�M[��ޖ*��ݚӣ�-�hCQO@��E�3~�uZ�EGH��2�Ɏ�yRhG��Oh�Œ6J�V�[�cY�T��S5��4t$���O
��H�J`�f�O��d�O��� n!�֫[�P�^��l�c$���Ie�D�99��y��J78Y� 3�BF��J ұ�S/��'f�=I
�+�.�rѪٍ!��87&�',���?��pb 9A�S�gy�O���(D`�y:&�J$KG�!C>�O���F/W�ͣ��Y�T2�@���i#���՞#<��3�?�+O��a�������F�l+�� ���e�ҭr�J�O&�D�O*������(p�"�Ot�SR���1���B�q�E$F���2�!#��H5�K�Z�ԙ�%��7�M�
H.;/tB���X���zA���nxC`Fŵ@��lk���O���$�rE��ɧ!�&|S��)��DGa{�)�	�~Ԥ��TcmaG�ɩ��`j�!"�	o��b��A3,��o��L�	��\���G�U��4��[-mR�񻁩���$�'�|��u��O,��ij������ɳ7����A��\]��&�O����ϖD��O�����,@e�-f���f���'�M����Lx:ypצ�%�8�c@�U�v �4��$�]a"�Ü��튰˔
�Z��>�6�~������MQ��8I��.D�G{��'V�k�n]*i�X,��꓍ D9��'����fC� }�≈�dF�yƨ���'�ҵI�M��\�	Fd�6k����'�Z��^�l��ģenІ�Ę�']�y7)[o�zA�T̖+	=���
�'b�b�(ˑE׎��#c�;��ȓ1�P,*���5�l�b�.ߡ2 ȓNWBeq�J �0X3��^�����B�v(��2d�I�7�06����ȓY�xp�A�LX �6w���ȓD���R*G(���vD��E��%�ȓe�t���X/2�d�bE�Z4�܆ȓWҐ�$�]�l�Z�	"�͌AS^0��Kg"��T��c�� 5N���<�ȓs5���T��Z��|��aq'��ȓ0)�Hb#ёZ���͓�9��ȓ0�����i.�Ej�Kj�ȓ*��P3r�CbPʉp�KQp�P��Fu����Z�#�h�i0^�S�t�ȓFܨ��n
����a��t��ȓ=� �0�o�	aܢ`q�푼}r9�ȓH7��� �Uzh�٢�Ϣh�h5��f�6����ܿ8�&�"��PL9*���d+biJa�Phz�xQ圶^����l�
�җ�B("�Y
�Ȕ�7(��ȓ
��`5�	%�*Tr�j�	�~-�ȓ�T�8��/V*~�GMRg U�ȓ 5��������1�^�88��n ��-ʅr}LYa��ޅG���ȓ ���r�	'�ԍ�sA�>a�j�ȓur���$����a���Ց�jՆȓH!`5�
�y�d @S%�[H����2{��Ru�f�D͐<fw�h3�Ǖ\�<	�P�5��iPc�L> �ySC"�}�<� ��Ag$�L$<t���X1I%�z�"O�B�l�O��"�c��N����G-# ǆ����j}b-�>����e\H!�EI�-�r����C�	
��ZE��2w��¤+ŞӪ��QA˫aX��j�GZ)Ȱ=�@N�q��Ic���+eD��UB�G��Qʔ�6���j���Mc��G
��Y�'́�&l���I�B�<��'ϴO�f`
�mI##���a"Zv�'�X�"[4}p�l���S*Y
�Zק�=90P�a��C_$�C�IdX� UL��4�" ��f�)�r�%"Ǘ�Ohy�3?� kAG���妋 ���c�O�<c`�uXmp��8�.�D@ 5�aw���Ω�A�'|��[�CX��h,#�hV;(x�zӓZ<�1����V�C�i�����lY���c��!�'>�)�"�9A� R7�S=#ۖ�S�y��R?'ӆ�g#ћF �"}j�ӱ��H�l95�*(��JP�<��M�b\2��0]�}���(��jF%B�+�	�@)`"|�'i\�Q&c¨��}�@[>^VX��'7v�c�HyX�E pKжO�P���cV8�T��%_���䛬\D�:7I�M֍Qb�Q�
�%G$I�F��Cq�Ż��i�pݲ$���V5��� F^v���'����1��.B�ܠ(c��7Ob�r�y���3Gr�2pX-�"}
@���B��9��a�
�|�<y��&b�nH�C�e�9�4L�St�Lb6�<l�I�=h�#|�'���/�tL!�� N��%�RLu8����J3�~�SRik7&Q�rR����h��q�吴rk�j�!$lO(�h�/w�֤Ч��?{8НQ���abC�ӂCپ1�W�R!5Sb�c�⟖u\�B�YJ��K�a�@�|p����~[8��%˻ V�"~�	��ؐC�e�F�X�%�cC�	 O�,���i���2�k\ ����-K�P�V�'X �e�=�j�h��ҽ6�p��I2���IC��<�C��Ѥ�DV�D��AQ�e�<�S��K�dt�����	 �Xc�0	P8+D��������Ht'�eŰ��pd\#AH
 �"Oxi!�B
�=��l�*{/Z�)���4���j$�|�|����qP�H�Cj���,D�$�̵b�BLzW��3!�<(��O�|k�)Ŧsmj��T�e=l���HH�6�&a��<?�{`Ro�s3O�Z� �g�ZܩrIۅK��2�"O�! 4-[�t�i2�(ՊRs�MX��d��c�0�h;�6��G�Bw&܄pI�_�T��(��W\*nX1U'�6-��������,������ż`�>�A@���%��1�oεu�!򤐟a>]h��:% 붭�8(*!�DǱ4���"j�|#��S��>Y!�d] ,$t]Q��Ċ�l���	4L�%��B�q�ZO�}��+���`�.�Rd�Y�7�_�~�����Z[ Qj�J��r(�}q��Ɏ}�p��	�R�dyj���=�'h�/H�rT�a�')��r�@r��X�rH�#����x%�a��g¬5TL�b3��5����aS,�2DI�3���6��3`��?Y���2ʶx�3�'K�ހ����ZB���P�"��U�*U��Ȥ{�X=����N�6	u�S�:Ԑl�'�>Q���Od8krl^+C(9+�.�5��T�8"��F�TD�M���3JӋp�
���*I>�?��<�$�H�1lO6�qF��4f�qj�#,��x[$�9���Gz��;�H��6�l� �H��|�y(We�;#��g"O���eXM:d������4V��߆$�լS�^L6m�fC�����1hAC�eV�i4<�!�6az2��Zpْ�;M�����oz���]c]3�E�N�q����:,��Ex�7�SI1��Y�C��05�,�A�c�4�$�1]��t�ؽ%�0u�$�<��?�x�bH�H^���q�ɼ,	�D'�����~��X*Pl�T���#�/�g��!��BE��BQ��{��s�g0}J~jJ6O�M�H/ �\�a�҄Y'ǈp����$E(}
� �̛�G@����s@M�
�Pp��|rH]�J2Pq�؜y�l�B �����'��0i��·2X�y�#Ժ}6�:"�dO�M(���O��b�>IǬ�u\csi������fF;hP�1;T�EvF�b�]�I�fc��"D\X̓��*bKA7(k,q�GP8)0,���I≀0�`�b6u���B17��'�AM5u���2��M1gx8%�x�ޙjazҫ�*4�:�	�M�&u��*�dX�	=��t����V�����S��ߤZ�D��pf��5L� (�.�'5{ʥ�"��]���I�Aݾ2���#aOҹi�|j4$��Z��ɫQaXh����p��y'(������t�jĠ#�V�!��'�q"�X�H����ȁa�y���5V!Ȁc�]0gB����푮��c?H=��Y�[/������=W�ɰv�űm~�t��Jț;���w-,,Oh`���ܲF0:�(�EЂCˆ����oH�,i �ө�,:��|��ҫ�1O�y�@ ɣ0oʰ��ĉ
*�������Px"˚2-�ZɚU��]H�: �]-n2�'��<���d�C>�xS��,+J��[U��V���n�=U�L��&LOXk3�Ҿj�&���Ί
䴸�
��%�>�Q���L���kp�$C�2v
�����
N���O�
3@�'���笚�%�|�(�-��7�$��y�%��ww%��銈?N�HY6ć�',�(��
6��ah���4$��ʙ�]͠aA%��vx���@Sr8� �͕.+V1�BZ�B犥1�G O��]�j���D*p�Hzx�P�0C�2_f.IQ �fr�� Uh<Q�
�$k*�J�(O�:��#�%/���'3R%ȗNP�N��ɹ$��pI0"hM8�yӆ�� �$��(P}؞p�*ã$�cL��0�(�MW��LX�'�44h�J>Y�/��4i�h��lPt�i��`�)�F��R`"�Du9S*�5r��>��NW�\;�!��Z�%lm��\I�MX�Y�R���>(�9X1�� U�F%�A��%h�h�*��UC�z­7a�T45�]%$k ��R�W�\jq�CU#�T@�P�jx���M�{�a�H�3��F�0A�1��,o
��I�'V�A1��{fޙbE�T�#݂���O̽1�R�p�j�/H�	�9�u	R۟��i�V)��K�6��d��'�2�Rf�(rf9������җ���^t��y���Ku^u�!o�3J�ȝc�D=��OI`V
Ԧ0Ql�Df�F�騰�ILJ��.��͓��]���I(+O"0gHF?F��*�d
��,���,�1d��eL��2ȦQ��'���%���a�g����'a���G�-3p@=!��F�A[Dێ�DL��&��r�T5 ,h�GlՃW��%J�h�<)^���7J��i�L�0�B�0CЁZE�s�l��V��U�'�qO���`��5��ݕe����&��bs��k` �(��$�kK8(�'��}n�@�C!
f2r�xr�O�<��O���f�N )�u��1T����!iڞ,� LK�Jx��т�.щgᑟd hJ�`ֲ��3�6	N=	3e�إ�E��;T
Y"&TP^R �b�\�X<<�b�B��-j�ؤ�A��{�
���ӡ.��|`&���D�F��m�<�����?eGЗqFh�p��@?q��+}2��&"F �"�V�sGʤ|sm �A���se�'#��rQo�Z	�MB��i|	]���pUg�!Z��L@��)���)Oh���3�~�y��6$�~���e�!��R�R!� �n�`P�1��c,��ğ�QD:�Ca,�p�8�ԢD�/�(���Ѝ �X1�%�^�ą�I ,�ܐS�,o��}�B!�>Q�U��E�b�:$�$քU-̓O:%� Ƥ���aL%�d�(r��T�D�����8�tD��F"�J�yrL���"�Hv"Z!�-��#��'�$d��cJ��*��M6nq�91@R(�p�2��ߌB��e�뉌F�}X�B�J̨�ף�L���j�i˧E�$)��Ȝ�9����dvD��$��{�Ĩp�E� o�B�9v��X�T�@�efF8)���>xp��P�%�F9+���G�p�aÀ&��C�NK�M�ϊ]����I<��Q�U��a��AӈeR����ѾHr�� #U�HG��sI>!'E�Ǥ�q%ʈlq� ��lܓW,Z���o�UH�LSw��=�i�=9`��^b4�`�*Į>[p�@�m�Z�	,g�ŔGKP7Z�d�2�^>-l�p"&�<84$r�-\&�=Y�mˠi������I)��
�%[����м~1�������a����'sqO���#!�L A���V0���9�y"�B�mB~a��(Ȅ~�恱�	W,M(E�*O���� OA�I�L�ga�� m>hR g�5:�Ā)ү#a|"\�>M�BP��_�8A"��U�<ݓ��F�$���BK�x�#IY��������#�Hő�B �I20f�Ĳ��7L��ق��*&���<a�aJ�M�aAQ.
�����~b�!?a�3#�p���2���)5�t�.�S��9E.�O�������hS�3e<A���ԝ���φ.��y����{G�����Y���To _[�H�$Gb�򰐑�N7�y�R�"9 u��iU�_���u��>� t+�@�9Vd���W\\����^k�� �-�ebȠJ�0���
�2 (�� O�,�a�/;��x���G�0�����U-5/��g��)�z5
�h��	�\�PǓ?
�+U�M�7��9C�$�?z%��Iv���H�����[�蟢o|ٱ#Á8���pl�A>eRq}H<I��T�g���4&��@C�B�<�+D�-ݨ�a2ECT��0�!}�<�V�
W"k�J�R�䄐���s�<��
F=!V���ҋ)�~i�׉�r�<$k:���,�V#��sѥ�D�<�"�� (�`�SJM{f-�p�\X�<�抺c�J�(��ɤ"+��iQ��_�<�0/D�D'ꘃ��K�pŠ��L[�<�c.M�
�D�I!�G�Z�*p�Bj�L�<�e˃jz�C0F[�Wj��9��E�<Q�ł�aX���!$�r!�� G�<i�OѸ���C��[t�b���D�<1�� �ވY�GT�0��r�+�I�<Ip!�i��I ���V9:`�H�<��eV#8�@Ļ ��U.f���'VA�<���I�|@�:���O������EC�<�Pfż"��<�Al�){
�Tb���|�<aM�/��QP�	f�|�q c�z�<���3���aʤ�.)�'et�<�tN�*H�(�B�  ;�p3B�]i�<a�B41I h��b1^��(��Ag�<��dɚ�(���L˪)tP�cw%	g�<�aUq%\�q���mb,X���m�<A��H@&�uq��
yxx����T�<Q��_$N�<CG��?��U̘O�<����%8{Xur!_�24�PBJ�<l8]`(���@�Y���DI�<�!��8f�$�#����y���B�m�<!Sʃ��a�Aɔ8A��N�<	�jD�nK��qՇǑ@Ab�P��K�<�n͸C;v���ȅ\6LM��%�a�<��O4j�e�����%��kWC�<Y�N�#?��SƠ�|���:V�Zw�<�f�l3�%��ŕk�q�A*Gp�<����
V�jl����ppbQ2��m�<�bbL�!|���C^�t������N�<���ȟP͐mi��J< |���%m�e�<Q�o�q�0Cc�
�hxyc^�<����P:�D�E&��y��8v��r�<�DCE#�څha�^��`d�o�<��N��g<� bgj_�D�ޔh!c�b�<)�i�&a����!�--���$	�a�<q�L�B��L���� ���P]�<�&���j3��3���Zp�EۢO�}�<D��Wb�A�"���X����;D�x�t%�-S��H�fk��<����e>D�t9��\�:���b҇�0�xpʧl>D�زS�ݣ
�p�h�,>=��@4�:D��8�&�e�&��A��4�-�aB8D�|��D�L)�!��+۸~��YJ�K3D�L3��K0�ꕆ'|o��:"B2D�xzSa��/*�����W��k�$&D�l
�� ���Bg��2���x�E D�`Zr*�8z��,�)$��IA=D��:��|���h�` �9�4��Dn'D���5�Ą��1ݢ�:M��&%D��
��S�~�KU�^d�R͸�j=D��k�!�"a�cæ7+>�9�E>D��+�$K� ��p	�6�T��`�'D�t�r �5�pk�$W`����$D�� ���#��rT6���cO�Zjh�A"O�m@r�ھ.��Y3���qP 	z�"Of�!VO7_(ԊP藥WS�*%"O�q�@4Z��5.��}dF�Ң"O�a(��H�j�X��u��YO��"OpHh��κg'~Q�s��k��� "Ȏs��äte^1��f=Tي�"Ob͊���f�I ���#�6�E"OP�[#K^�`;�}�����+�\]�b"O�m�`Ǎdh~��#�����Ed"O2�+C�ӭ8��Ȋ�AU>"KPqt"OX1��c@�g,��f
+N.�ͱ'"OP=�%I��m������=B<���"O�2Pl܌H�(����A�h$�-{�"O��A$�(/?�<y%'O:QdD�3"O�A*��snv�S�e�.��a
"O*LPH��O������v�.���"O|m�@���(:D�1Wd�g,-��"OΨ�4�֦X;��sb#E�#�Dت�"O9���&KӬ�0��Q(p�}���'Qў��@&U4P�fiP�C��G@����0D��I�@K$�x�I������ǂ4D�T� ��n/��"%�/un��g�&D�`H�+�=��,�Q�8`����M#D�4���5�<٢ud����q� D��B�!N�(��K$Ԍ|���
!D�|�ACA�>�A��^�U�ԶA $D�l�%��&q�^Ṥ�X�G�d7j!O�#=��j��aQ2�#])p�x�&_}�<a��S6>Ύ]0��Y�D�E��Rq�<Y��$��<�pJ]%��Ňp�<i'� �:�>mA�R�m���B�-�m�<��b�75k�i���s@����Cl�<9ul�?3�Ρ�TN0\@Pt�f�<Y��;+�l�d�Eq�Q	W��c�<���$A������'z� �dv�<a�b�ibx����w��0�f�r�<aQ"��~I�4�MmĆՙb�S�<i4"^�7��	0c�
��$`���c�<YQ@O)G}�d��T�2�BY�'��^�<Q�n�S�$D��1q�V�<����4�F�zA�M�"N���PK�<y���^���E
�r���F�`�<�`�d?� ����^�p/$j���.6蘰�0U�l��#j�T�Ɛ�ȓ0eHx�Х y�����%��\�ȓz
�9"rO�<�L�;\|���=D��J�! �#ޖQcOt��E�'D�p���	X9��$Mh[�y{��!D�p�����[��g�L�+� $ʤ�-D����]3Y��)�M��NYJa�7D���'�0�ش{d��A�Ů8D�8�� �Дa����z�� b�:D�P�t	�/�(pٳ���&�P�7D��*�n�LZd��f�3b�Zy:F�5D����c&������G�R���)2D��b� ��|�3��-6A�`�$D��I�>p���H���Ci%D���A�.?���%#�"��t`l D�`z£ɮ$�8�Q��[�xF�1D��ڃǕ�B��ã�<�r�p� /D� 1@cď	�|���̖H3`���,D����Eۻ08 )��I\K��0�*꓅ȟ�2G»C(�� r@*܁w"O� �xrэտYJ���E1;0d���"O@(l%+��ԑu
��Y��4I�"O�kr���B�o����"O4hi��._�Tp�(	�0�`B"OL��"LV���������r"O���p���[�>`���H|z��"OY�G�ɱf���>h�a¤��8E{���A<w^н[䪒�������̩-<!����>Ϛ%[�Əg]��� )� +!�
�A\z7�TFS�XT_�^u!�$U.,��K$+ LNt)����!�ā�D��T#�J�f�֙�s�@W[!�$˸8h�i5oN�X��fގ/W!�d}e��`�r���/k
�`�"Or`�B��,Eǌ�� ��L�0�u"O(��$@���э�/#�� Sd"O����DL����7�1�Ru�"O�u��EF��<���8�i)4"O�h�P�H���qE�={ ���d1lO%s#AF���xd#�Q��-Z�'�剧�0|!��M�|,0,�)ռt4C����P�t)��G����҆:��B�	�a�Ih�i��}��%ҥ)�C�	�`�\<q&h�	вA�Bu~rC�"�]:w�ޒ!�>�"!�N�&�*C��+l |����f���cD�0� C�Ɂb����W�Q���H�g���B�	���)Ձ[�Q��	�K|�B�	8	_l���ݍ#���yf#�y�B�I�B\�����FP�� BĨ�~C䉎"����$��U@@��(A�:�^C�ɂ�ΰ ��^8���ƌJ��C�	�d�B���ğ�̀[t�	�-�zC�I3_\M���<A��4������C�xx4�ʖD�.r�q�g1,�B䉘"�,�"lG�5���a��+P4B�	)&ǦYc��RdP]HъLS�B�	�Z�B��3�ϓ?�(Q����B�	�SY�t��B1\��4 ��H6&�B�ɶL�z�ɖJ�(��NF:�B�	5�^5��$�ÀL2c�E�HC�I!]֐�[3��?�*Ⴂ��B�DOt���/�FIh���^%L��w"��"��~⠧��)���w:TA�rx�ǆ"D�耰
K(��f�Õ�����<D��@#
�3%N�Q��&)hv��+=D�;'F�=[��rѪĔ(�1qE/;D��ѕU:XX�:�`>��t!%?D��o�IX�ܺ�@�Q=t�z�"D�(��H��\T *��S����/>D����%R8x�Z��<T��i��=D�L�5��0��� 5�X�z6�hO8D���@�+�� :�fĨL|$�A�6D� ��Ԫ5Ѐ��A�MJ� ��4D�<��-��Z1�ą=2�F�I��0D��J�/�$}Ј�Yf��5Jx����,*D�$I�IB.9���{3�ӆ�J�P�@)D�,K��Uitl�K娔�vY��Y �%D�t���W�G庴�өǶ]�n(�'m$D�p� FM�1vf�"uDƐI��4��"D�$�_8����I�-�n`�`� D�@
@@��p��I�ƈ>�T���?D�Lg�*�H�����6C,xX��=D�dzU�Y]_= �C
j��\�R�9D�� ~Ua�ćP $����c]\�"O�������kC`	��-߂��"O��"�U"z��0�J0(5|���"O�8�C�L-�|���%j(Ƞ��"O|�Q㕴��@ ֋G�qX�"Op��S8u(Ѡ��$<�L1h3"OʅPA�Թ�۴�IP�0��"O�Ź�� �N�UIP�D�!�rY*""OƐ�ԍ�,WHd��#Gۢ(Q�"OLm����"o/l$���x����E"O
���O$F�X�)�c��=��[c"O\�%��9(S���w��#(���"O��ȡeX!�xy DrU�f"O���D�F3_W4$�cȕ�$�*y"OV���
Ji7��@1�%7ox�۔"O0�1���y�� Z5*æ��"O�5�Q�jj�#g)R�G�dx�'"OXl`@��=4�dL��N�.��� "OJy��A��@$��⤇L$j���i�"ObM$Gζe
L\��&��T],c1"O�����E *(��2�I@����"O�L�P{ ���w56H)Q"Or]iH�	�m*��[�B��@(w"O�,�� ʒO��$�X ��H� "OJ<�Db+�A�EW��
�"O��)��#*0��e���X�q�"O@�1�ڢ�Ҡ�)X���C"O��V��XRF.EZH�M�y�ֈK92QbG�2y:�	q�2�y2��}^tHw��'p̒��p����y��[�KF���kʄn�p��D��2�y�.I+(�R�+f{|��D%H��y�N�z����
3W��S��G�yBJ�	&)H�c�L�<�2��y2�Ӄ-s��
(֕K,@CR�
��y�	̘;��]�f�E8L�U���R��yrl�^�r[��L)Ll�"�+�(�y�~��-pD
�|��!B�@9�yLеF�����F�zX�=�@�V �yb$��U�b�Q��Y��Z1��A
��y�S�.�8�ȑ�Q!v�nE�4,��yr�љG2j� �C��^�X�U��y2��~�{�(��.�Fa�dΞ��y�i�$z��A
bư� ct���y���9SL����C���(j�-�yr� ��P%�@P!-��h3NR��y��$5I���&H F����>�y�l��w��dc�鎪4B��n���yB��L�R�F!?��S�FU��y��ʘ�e�P(�:�2��@.U��ybN� n��5��`���2�M��y���U��!3�O%
d0�q'O��y�ם�������v�0](p���y"Ɗ+�@퀱(�2>5\d������y���48���%Z/9����ƞ��yRJ՞^����'�$S�x���;�yRb{@����H�1(^�e"��,�yr�P$5��1��ҧ%l}��-V�y��3GP,�r�
>����ۊ�yR��j�1 ����A�!Y��y�F�#Q�T��JΗ�2��!(L�y��B�	��ٲ�ɣR�Z᠀0�y�).\��G�^tp;k�y��BH�\Z�@ےY�x;��>�y
� 
q;p�ȓH�bM� E�(f�z��1"Op��i�R�Ш5c�80���"O��Bsđ.'���z�Т1��p7"O^-s'rtt	Ӵ�M�1�4�I�"O������s1@�{��\6MhI�"O�!�̋Z�MJWo 7뜱c�"O������3r��1 d�f\8�"O�����	2�ŮZj����"O`$	r���;�.h11Ú*fW�|�6"O� �b +B���1k�"'�c�"O����I�X����!*�0.����"O�U���wJ���hY4cbZr"Oڜa�e�5&��sG'$C�A�"O,�/M�8�Ǉ��;'@��@"O�e�i��Eixus&W�1K�"O]X�	RR`z�H�ٖi���"OD�p�L�V���� �DZ*�;�"O���W�X��
.�E�3��<�y��հj?�DJc ^4:Ҧ��y��4 �@5�E�5� xA$���yr�(mh��$%�!
��ӓ�y҈TG*��h����b[��y2H�1^�D����[�hհ�k&��y�$D����c쳒����y�M�+M��㍚�b����bJB䉗Z��d(�Y�QRT!�'E�gw:B䉻d{:�	��I�[�ޙ䩂�8NB䉲d�0BM<��}b�^��bC�If�H<2͆J.�U� C��cC��"��0�&-C@X���>�RC�	YtIr�қC�v`���*M�lB�I9��a�!�3gـ=��>5�hB�='~�{ EI�-�h%��D�frrB��,W���s�6j������(hB�	80Y�:�6Ns.�#���%!3LB�	&���0S��w6Ԉ���ΥWq�C䉶3-��+ҭ{���&g� b��C�	�0,xAB��G����yg�K�]f�C�I�9�ba#C��''��BV���3�jC�Iz8����Ͼl�e�ǉL��fC䉇q�.i��
�G��m��∘�>C��	W�8{w�:X3�u#��0[�XC�	�9N��G���NaPꆉ~�(C�	�%�,s��+�N=��k�'G�C��>p<�r�E'm��Y�Bb���C�	�hS��E��=L���6��K�B�Hۂ�q%�����"�ǛX��B�	!ez�qQHJ�a;�LEjH��B��<h�JЩQS�C�nL"G,� @�C�I�I��tQ�"�-mY��$ńq�C�	�  ��L9V��|�����C䉍s����/�Wol|qV�Y,��C�	Nk��EWdy4([s�يO�BC�	�T��A�cl�@ҭQ0C�C�a�~e	G(Q�� �Q��n�B�	�[5@P�U�\0`�������U��B�	��E�*U�1<�����B�Io]xQ�i��&(� �Gy��B�ɗvK�m�7�@���E��$H��B�I�hܑh�z��B7�W4j��B䉼"�и�F�%uA6��5��q�B��5fn����-�Lp���Q���$U�s��L��T�8X�&M!�	Qw�Q��6V�^�:�'լ;3!�� �� ��Bc�@�rhF.m�H��"O�L��$BI�&�i@�_l�����"O�p�4y�Z��2
I�dEȼ
u*O��BW([�E�� 孛�P.J��	�'	<�Z�nT�N��m�$�A�O8AR	�'��X��^��48���oX����'�p*�LG�Px���Ӡ�a��	�'x�ti�m*	tM[����M	�'�TZ�&_�	+>H8	�� $H�	�'�0D����m� J���%�. �	�'��(�Bd��'e����d�-'�h-a	�'Ă��&&
2<�.����ڡ�5��'[F��K�9?������Q4t��b	�'�*�jw��>�V͙��x@��'���ъ8V�,L
#��&˜���'��1�5�.�*-)B���|x��I�'�Qs5�� ��y9�Q�"�����'O��a��yUĔ(H�-�Q a"O����悑��󇘆O z���"O�8�����e�&L)Z�z�"O∑��;h=�$�1EK���yI�2V^(P��"E�F���͉��yrC�K�fi����_�\�X1"��y���s<�h1*'�������y⥃�܄�Z7O�	��e���yf	��7��6��FA��y�F\�kN��q%[�Y��0C��&�y"!��x;� ���7������yĕ�M�Ja�1D�x։� ����yrG��,npqgD~`�4���߳�yE�5I&"@�jNs8ب��lE�y2HI�p�PJ�qF����y"��8m
�KcB�F�@Z��yr+ �F��I�6.���$"ЋE)�yrFВu8�[���6<�JG@��y�,$q���o�0���顩ˁ�y�(��Z|%�9��:AC��yr�ހa�H��a��#>���F��y" J>;�$�a��N�r�Vi����y�'�|�АR�k�#z�lrDg��y�(��M�΀x�Ën��#�L��yr.P�2
n�Xu�e�ܘ���E.�y��'�аC/ǍV^1��'ݽ�y��qT.�J2;V�R���*�y��2Q/����M;A�\8�A@8�?����<��d\2��-"���4+0t�g���!�d��m%��#L	�1-�X����BD!�Ďբ�)��͹�<��!2!�Ą82�Ѫ����>�#��<�!�d5/N����S۪���M)(	!��B�VlaK��
:z%{�D@`�!�d��q;��*�
<������9��O��d<�61ҨЇ#�5��� �͏�'�3��x�/P%b���D�.y���,��y��N-��YW�#q�̱�"��yBeŚ!X�`RM�=n�t\���ē�y�c�g��iȖ/T�t�TqCE*�;�y2�R������Ⴤw�tYx���y�lɷa �<Ip�E{�p��(��?��r��ٟ`�.Lv'�uX6.3"�p��4�����	Q��xB�o8�v�`qn�* �>���'D�HK��]�x�xm��XY�xx��2D��k��N�
2�E�$�Uw2���%D��A7�[�_�<�B�#�h��! �$D�� n@�$)M 36�@�P��"� =��"Ob��$��40�.YFƁ:48e�r���O�㟔���<qS�� aTuˢ*�t+�i��b�e�<�t�Y�k�>����?q<�ST+�V�<���00H�|��#B��$Ðf�P�<�"�Z	lczL��ڍ� ���C�<��ϊ
`�<2�W�bӄLPJj�<����
��$� PB5Pc�ON�<)�"M�D"�kQ��<p�6�YJ�'Za��/(��Rj^/-�v�b%i���yB�[�ztج#�/R)�fD��a���hO���)ۭ>b�1"�8Y�-�"�B	J��{��dʃ��@R)����Z�\$d�!�5tlV�S�͌�-�p廒e ��!�I�N����!�U�9g%D d!���,J�����*s�r@3�b�cS!�
]~�4!�P�(bqW�P!��B1(p^ r�Oŀ ��DA��S:!�/UkDb�Y�A�fX{��2�y"P���'�p(y�,R&$^��f�$y�B	�'��d2�j�*�"�rM�8d��\��'���F��L�v�k� ٓ_ʖE�'�fHBhM��Z9��M)$��	�	�'���� �O"�#!�#��a�	�'�R�R��IM�|�ρ�L���ȓU<��
���;B���[&lԑ"�%��	{̓vqD��2��R�u�D,�	u�����<4�lֺ7Ezu�bf[H��<�ȓ�Z�31
�)N�LE�����L��ȓ��as���@ԋ��Ef8��>J:lҌN�o��B���,Vq��/#�����a��h�яK�-�ȓ(U�a���gD���]<W�:��?���d0?q�+�V�6q�cscʅ8��RD�<yw�9.K�X[�UQ�I��F�@�<	Y�&�*`��>\�@�$b`ŕ��'Qj,�p��:*��Y��-S!�Aq�<1�ǃ�tn��`�[�f@��Z�8E{��I�E���3C� _Ζ��a�T�B�I�8UH��̶���u0Wb�O<�D'LO~�!@���@d�h �-!p��"OLaACM&��Y�V�P�"O0��S��z�d��5F߫7�V�S�"O�X����(Q��|q�&\�>jF�B���t>�Ҁ؆��и���%m��C��/D�$z7�C+,u� ;h�5t�L�R�*D�P�bW ]#Zt�h$GʨC���<�����(��1+c�>+�=! hZ�$��}R�"O��JW�щT?�����H !�H�f"Olek��GX���r DA8=��9*�"O ,�50g�#WA�x���;�'����v��.��[	K�^�p�"!D�p��Gӄ
�R�;��?Vz4	�w'=D�T���i���a ��uR���O�=�O�1O��[�P�:m�����YDp�z"OE� �= RD�q�qC����"O��(� 73��Y3g�/.;��KV��Ryr��H�T�ȡ����¸Z���!�� %Q�b Q�eL�2Rny6�I�F}!�E�7!UJĮ�>�Sܗ��u�<	��;]?vE��]�A=b�c'��lyr�)�'�N샐��88ʖ��u�L�o�:��ȓ����cN��(���6g����ȓ_��Yf�G�?"0��a��6��E{R�0D�� $0R��ϯ���f����%"Ol���A'8a�$"�_�����"O�����;�􍳣"�%D�:�p#"O�U#� "H���7�HnA��H��|B�)�� k}K_?�p< T1����"O�yؕo؇)`d�ه�@=6��l�"OrT8΀�w���`�bu r"O�����#*��T{Ť��<��	[�"Oz�zCH)"<>� �� O��a!"O@�Qlz���Ç�M��"OF��g�ս@�h$�fh�n�$ ��"O���$�D�y�NPK�!�i�B�j�"O�p�C"����{£D
9-M!�"O8�C�=!����V�ܤ~�t�b"O6@Q.m�|���߅+	$U*&"O�Q�iU�bcBm3��$�j�R�"OfAs���1Y�pYj�b6�<ua��i>�� �i�Z,�Ӈ8���PU�5D�$#���K{���f��mӶL�#.D�xi�f�?|t���� *(j�,�./D���F��1F���N�5�����.D�0�4�Y�Ъ\1b�[��vJ/D�HC�kE14h��`$
��p ش2D�|Pū��B�~=���ʴcDB�KP`0�	N���ӎX�(a�d��.��ġ5�9��B��<j�9P�#���2J�{��B�I"u��y��o#qr�%(S��B�	�U#� �R��:��(w�^��B�ɾu��8(�#̌o�T�0Պ['6�H����O�Qq`��@�HR$�Nc��ՁDk&D�$	� �&n=��Q�l�<���{�e�OL�$�O6�=�}Ҧ��?;�Ι1�K�W�09cgHnx���'�M@���t���v�?cz�AH�'A�yJ0��%L����6JRo�. ��'YYs厉q������{�b$��'���#�d��� ��Q"D��'H~�z1M�;� ��b)���H@��')��P��ȺD| q�CZFX���'C"�I]�'���1���%&ȡP  $pVͫ
�'�l)�@Aכ%IF��UƐ2c��*
�'|����X�w"��G@A�P��yC�'u�epG���0���9:���i�'����RHZ���։.LL �'��A����u	ģ��!��hy�'����#\�5�R��f���
-���?9��0>A�ʀ6��z��2t*^<��
�W�<��)@4'J�JB  ���t�&�T�<�a/�$��[5H/U	,��TG[W�<��e]�X+�(�����.}����m�<�d��$�&X8�
I�u{�l�`$���������%h��7�n8�&1ړ�0|ʂ  $/��uKS;(��H�^yb�'4xQA�s��̰%�H����TV��#�Tr�*b��"y��р�;"O��Mm����*ăb����
ġ�k�+s�\`�2k?c�n��ȓ�R���P�A-��ѓi=��IG{�O#��2�:j<LqBM�5�@!���x�-d�VtCG�K���5 ,�&�y2���2[Y8�Q�+蘔 6N���y�#+ߪ�
��;2^$��*��yB(��F"��Α�+���ӴG��y�Å�N8|�͂�!��*��-�y�*X�7���yw� ���YX�l��䓇?Q���� Du��(Z�.CV8P��;��PhEV�����+�q�����!�k�4��B䉭D���s��%^H�炐h�B�I�F�n�@�%���jvOM	q�vB�	�9c��+f0��i)�h"=�dB䉊d� �^���r!I���B�I�]�>U���%x:����4�S�4�'^�	�@?�\����
�x�Rd͚�*�B�I+@y�t�p%	�J^���خ�B�ɾ}���@�ێ N��zd�jxnB�	$yK8�SSZP��єƂ�5�VB��3|m��k�צg��L�2��V�:B�I�?(�#���y���ZČB	K� B�9!�d#&H��a_H��ɜ_�C�	�)]�ɂ%�؋(,���b��/��C�I�����RnB�7k��3W!��8h�C�	��<�Qq��{0�QbHII�XB�	$x�P*$ȈIҊ�Ȕbűr�.B�ɃR~  ��Z�!���&��B��nטp��E=t��ip��3!s�B�ɔC.��E_�+*�aI�4|0�O\���OD��	¢��Q�F	z��b"JU9Bb!�P�S�Jlڱh�2��B�Z!{2!�$U�;��ɚe+��?JY����D/ў���&
؉�!b$>����%hHB�	�PB2T��I�U4 ���,)�B�ɪ��! -�eSra{r�7Y� B�	%nJ�yK���Yİ!��-��Orʓ�0|����`�2�jG���L+�F`�<ѱ�Ĩsn����^A�e�UR�<1Ů֑Yk
1K�	N�j��5Ay�'���S�"颴�E�+b~����C�	'�R�%�^�,ЙSo]9f$B䉛?U�����İ �>��d̆�>� B�()1���F/O�eLD��A%Ħw���D{J?]Y 2�t�S� ��J�*�N�O�B��,mܮ%�����<��	�/�;�nB䉉N���I= ��A�q�ۮM�?���	5tE�T�2m��Iޚ��,R�z!�D�dі]Z��!Ӯ�#�'t�!�dєd���p����������X&]!��kێ�(�CK $�F�@�����O^�=���9��Ջe"��GN�sk�m�1�'�!����C~ ����0o����G�@f�{��'���0q�l�W��>d[��s%-�'XhB�	;`)~A�V�K�,�qC���>f��C䉾q� i�*N�'^BM�}1LD��'F����=�|�n�{ *IR�'�
�S�Z�"M�l\\���?�h��H�����F�s#fĂv�ŝ�y"ğ�`�t�i	�dǂ�j�D��=*O��	�*q�J�'��d=Ƒ��cW�Q�:B�		PZ�4�r���uv�y����+��B�*���d 2&�%�a��"rFC� !�D��C0IcX��2�ǅ"�C��m�aa�a��s�X=ˤ��+�B䉁[����R|��Ŧ/�nB�ɷ|^�x���O�(���KF?@ʤ����O|��{���X(M���Z!nϿ#�
a��+D��1C�S&�r$�	c��i�m*D�h+0OИy� 1����(�[�+D�L����.(Mh�n�#:���4D�؁��B�E��|A5 ʉ;�h&�$D��R�͍�,�vM�D$��D�,�1F"D�� ��IĈH�<�t�p�ɒӰuC&"O��V�
% ���s�Eƚ?:�ؠ"O�A:6�H;:G�HaQ�� }4Ĉq"O޽�'�tH�3��ϐR)���"O����jO�?o�!����"
XLc�"O&x:�P dy�hIV$I>��"OT�Yһ#�x�D�kL��s�"OD�yeB�]�~1�ƏG�&��)+a"O.�y�E�5&j�:�_�ĕs4"OF H�A� ��q�aM>E�Nm�f"O��qenA(���bMS�\��"O����aη/ފ����H����p"O�!0��l�@q��`���P��"O^PU�,W_��G
N�CE"ON5�,��l����p��,�db
�' H�q�*�8B��	���Z�k<�3
�'��5�&	ں}-�uc�J��4����'v��s���fL㤈X�#YF�A
�';LQ�FfӒc��Q/ƪ!��+�'�"�Ç�9e��*�e�Y��
�'�`��@��2"�"�!1�
�� j�'6�y��ڶh��c������h�'P�]�r�l�L|ӧD�vcJ)c
�'^,�Q&��p5H����AܒM
�'NZ�;Pģ��'��8)K���
�'���րK����b��iU���
�'긐�FD
J�R}�
��vr�{�'�%���y��dj�$��x����'������?9̦�2&��jk��	�'��� G�Ǐq���� `)�����'��r�*2^0��(��l�ԬZ	�'Vuq2+�?� I��>5�L�	�'52�B�"�����R��#\O$���'; 5�p�@x",�'[��9	�'W ���U�pC&D��hKlȨ	�'�J��RN:�ʠ�@�g��|
	�'�HC�0F�$�q$�+u��K�'��L��C�5}�
&�гo%���'�v�	� U8 5�]Ң��&�u��'.�5���1�-a�O�����
�'���2��y�@H*¡��+��
�'6 �S*_ r�0[RD�8�Lq��'�h�kE%�����M�@�-r�'4�x ��׼b���W�ִ_z���B�'�F��5�L�%$@�#G��:���'�d {p��'�F�AV*���'�7K�V#�Њ���'�Pi����$&^X5h�.J㪵��'�h\Q�S�W��� �9:���p�'5��Ņ+ń�*uN\?5�`��'5��mO�0Ԉ�S6$Q�ݨ���,O�u�l�7s,�H���9-���{3"Ox8��FIqJ�dD�[�>���"O4�� BD��+��.����"O �j��S�#L"�p�j2F^���"O�d2�# H�b�JRE��+U"OL݀����)��a�I۞N��!"O��i퀚 �8���J
hl���"O~0�@ˬ�`�N�Pej��"O��b�*B�^��"T6'tE�@"OL0f��Z��Y� �D�ָ�q"O�8���F*a�wm�7g� d�"O�"ckU�q�P%p�kR�2ɣ�"O��XGFD޽+�R�\%>5Zt"O� 8$9�"�6p�ƙ�p���c�61�"O��Ҍ�it����9�>Qv"O*�s�\ ێCa�Ң\}���"Oh@ZSl˾AS�=�#��$Q�4"O�T!� �i@x٨��N�=Ib"O.\� ����~�b�&�8O����"O��@�cƠ�~�9v�j���"O���5�&?"l��S� f���e"O����@��bFHU�n@�4"On��0�D	~�d��DbݢtN�۔"O���4���4���łF�~a$�"O�l� +Y�R\��pr�TDY>���"O����!Q�� D`�.Vp*2"O(��2��l&��Z&*�I�=���'F���3.R����[5�T�0���!����|�Bт�:���K��	�{�!�D8x��j�ֺm,��y��s�!�9}{��
��c&ѳc������GiD �J�?<�4!c�	 n�BC�<_����C$�љ­�b��C�I~��r%W��X�����,��d�O��D��Y��k6�TA���W��RwC�I<f��8����5��4"􍔟	'6C�IE>z\`�(ELXL��Vj�6��B�I.�B:R���>�ue:w��B䉌\o:X�\�;/2(i``��8�NB�	6�H3���'>� ���JvC�I�&ֹ:��A	|���Ƞ��"<:�B�ɇ�����t��B$Ǭq��B�ɇ�\DB��A�^Pw$
 [�pB�I @�0bA&���t#��@,C�	$�$�� �A_�|�瓵e��B䉤Y΂((��aw�,ۢސk7B䉩lI�i9���(*\�	J��4��\��ɿ�AG/�̑���ו&�6C�	B�y��%�
�Z�V0��B�	�!�<�6%� |�`��_�.GC�	5Q����f 'Z��aj���&'�NB�	658 0t�ͲV�z-�gΛ# �B䉄�P���jN��T���U!�B�	�m ��TI�բ]�æB�	?�xmS̓�>��.��8�g�&D���q�B�U:m�.�K�����1D�d�d/�;�ɓFV:)N����.D�Xxr��%U޶8@�(�f��c:D��ծF
�����KT?��Lҧ�2D��y�L>��i�ǌ;`�ְ�'&	���B����-Cc�
��"aż�t�a��?ɏy��<�����1�L�ᣈ4
�F4+Ŭǋ]B�C�I�B�-�r�7J�<�WfC�^بC�0^�G-\�ؤ9�F\�g��C�	�m��q��-ä�x�Fꄅ.�RC��3u�p*��[�$�����J\hC�I��L�(
��S�8Ec�LC�ɇ]��H�&C�^���
i�/\`���O��@E|2TQ/0����1{X�J�����y��W�iS�S���ojuiq���yB���*�j��N騅l0_(�ȓ~��Ӕ!O�,���Ԭ;�zp��#�ĸ�+ƎZ ��,�2D(���Ɠ8RT�:L�O�B%�FYI$��
�'��H����mhr�Bf`܁I�~@��'Ŭ��N� b�h(�u�';���(	�'�Йxd��-�l8�����6�,@Y��� Ҽ�E&S�Cb��Ȓ�E�4nx���"O4�Lŧs<ܙsGӁ  �"OJP�c�C�W�L�#��&�
�s7"O�U�e�~�j�����L�@��d"O���F��V}ɖ��z��2"O�0�Y�I-��R�K� ��"Ozu����^T|1#"���+�"O���E�H	�xrS!�-�t4"O����M(�F��t��)�"OPA;�C r
\2�ͪE�q�u"O��Җ�AXE )���1LX�"O^�yg`�h�j,�2�
�W�b�"O6ը1j4���y�#�iT\�q"Oviag4r�F���7T�h�"Or���qcD���eF�1V�Y'"O��Ҧ��"	���<q�,0""O����冐"�b��a��O���"O.L�Ë?p�#!�ԭ�xظ�"OD����5﶑�PDY=>���C�"O=�4!E�5IMX�!% �4d#!"O��`���\8A�jN
C��k�"O�HRU���J%3�Ʉ*#`�PQ"Ot�Se!]�W2���(T�]�"OR<9��v�}�&�S]
��ba)D�8�fG3����RF0.��lZҊ%D��9�O� =F�S�o�pӐ���"D��Q	S�v��$"t哩bz`i&�.D��8��I;�t�:#�4LjD�R�.D���)�&<���uFCa��¦�1D���2���G��o�x�B�AF'5D���H ��Q����/�Xm�b1D�䁗�ԍ|���R%D��j��<��4D�4S���I�����[�긨��0D�xQ"Ɏ1X�T�6�š0������/D�@vg�}Ҁ�֮��*he8D�|�p�;H��l�tOV�RƐI�	1D�\��NL�,�Yc0�Ӷ�T�<D�l�R�=gb 5�Ñ�DnZIh:D��Pa�Ǣ/�V�c�+S7,8�k� %D�8��ꓹU����� 6:hKp/D�г7g�$R�4l��ϩhy���,D��b�d�O��#@�P�r�*0D+D�0�Roӌ���ƀX�1J
+D����S5$�\ѫ��]�!�>4z�n>D��R�U<�\�'�5"�JP"*D�x���3��E&�1c��O��=E�T�]�	p ���@� |��(�+߶,�!�$��W�"�����B�(�+@	�!��P�͸t"��D=�.	8���!�d
)���%s��<�V���0�!�$Uj�9��m	�3&�K6c�"�!�$�I/�щr'�1o���p��@!��މ��Q"Љ�
,�U酰��ͅȓT@m��Ӂ��`�a�׺Tq�Մ�W������(H,����燴`�-�ȓKdʵ���He���MH3N6d���oW@��e
�%{J=j`o�T�t��ȓ4:<kc��-94�!"�U�E9V��7o�	��fӣP#���hZ�ӐE����UK�f؝~ĩ�#��}�	�ȓYF̨&h�;�`|�Kևo�ʡ��^(��w�� Y1�81S��b�ńȓ[%�L C�V�x‹� -���ȓ�ZU'Wn���S�Y�yw�ͅ�S�? L�0���k��*�E�>#]�T"O�<�'�3@���dk��y��"O���I����L��w���"�"Oh)����"W�d���*��)�"OF�+aBֹvq:��Qi^ M���""O�DX���0u,@KƇ �R�@��"O2u�G�M#67����I	 �6Qb�"OL�r�L�Tʠ�cV�O>���S6"O�]J ϨV[v(IGQ'-���"OH������è(}���CA"O~%r���WMR�HD(m�f�aS"O����@�Lp�SQjN�p���E"OJXS�/X�8���Hԑ a��¢"O y��Ŵh�=��GӹQKL;�"O���Ol���EO 8�9��"O��(pE��f�j(9t%ʐ\2�刐"O(8�]bL��J��T�t�i'"O��x�(n�9��	O0t+ "O|����\#Z�4�2 �["<h�"O&�RGǿT��0��hS.g��z�"O��bD�тc�T[���|�؋c"O���Q�ֳK����å;h�R�д"O.a����\�5'Av_���A"O��K��Lh�}�l
�b��R"O*�� l�pd�y�l�$ߎ X�"O��A��;2^��H���?]�|���"O��B�Է]�v��s�x��#�"O�8c"�0}��-h�gڃ0�J�j�"O��c�
W�v����&G�G�*�+t"OU!�D�3�����*@s��Yc"OZ�wl[!\Ll�"䙊c:f���"O���Y�\���cDL�
U:��"OF1�0�̬'BX�A����G!��"OV���4J��:�#U�A�ӵ"O�-wQ�F�UD�R���k�"O4l3JX��XI���R>o3���"O���d�,H���!L2�0�S"O��#J�	#6U�5�=ʰ!B4"O������B����&�Z��vH��"Oʅسl��/pؙR\�"�;�"OlX�GjI�������*Zn@4��"O%�V��6���[�`�#m�$��"O&����ر7O0�K�o 5_�0
�"O��Be�Ւn{F5��^�aL���G"OD�	�ď.W_^$��n��C,���V"OH}�	р#�>����(�Ȃ�"O�-���3�X��`K�h�PD��"O���)��E���� 7n�p���"O�D�UF	 ��3a�H�$"O8h�� ��,��㤐�Lz��3�"O�����I=.h�ـ�P=?qL
j!�d�����M?^d���fqf!�9�"H��M��t1�ԵZ�!�dZ�}�~H)�]5�����r�!�E � �+�ǐ�i~�4R�!E%1�!�dQ1��!��ܛ%���v H(x!��L*:�-�I¾W�ȕ:'�#a!��J�2�R��!HO�m�lL�u.F_!����+}�i��JJ�����n�<OL!�d�%,���I::ܬPQNP�T!� 9�&M����L������
!�F�s��\ڴN�),y��-��:"!��( D�
5�N�5 ���)!��E�y(_�}����e��u_!�� �	�!&a������M�N���"OJ���D_==^�س�
M��`	"O�m(��)�@Y=5ڮE��"Od50��Fp��ꀀ����]0q"O�|�������#�d��=98�q*O�ɐ�#�m�N���*N�AG�0z�';�I0�
O�t2q"H)@�����'h�1h�C��k��Q�GO33:t��'�̈��C�76h@�'o�XL�8��'naE�B��*\InP�'B�
#�'9x�:�lY.X��h��'�0�Eˎ�Bޜ*��B+I�XY�'��<8f�� P��m�N��E��%I�'IÃ
��Д�J:�T)`�'�f�B1!V�`h� �S7A�� 
�'�(��N8�"U�%j�!`�Pp�	�'�4#���9���٤!@�W�	[
�'%�!q�'�xӦ99�Ǚ*u�y	�'���*ӬߌJ�*�(CM�!y�]�	�'�^����jd�
S���_H�R	�'I�%I�⎽>ؠ��ǂ���Y	�'$8LB&��H����ك�6!;
�'2���V=p/�M#��S9� 1
�'�*9���G5��b0�D�f�^P��3�- �A�kXԱK��Їf��� $×�ƒ fq��.G�2���ȓ}.ɑ�/� .@����]2u�,�ȓG�(����I2x�0���!|P0J��5x���U-�#7MDX��9�P�0�Ε!C�|P4���{S2��B'�`b���q�� ���x�0��\����S�P,SFV�Uf<���|��t4Y�� :4l0�I����yG�(.��8��e�3;�h"����y�[6PԊ��X�}�6`A�/���y�$�8A�	y�K��z��C�J<�y�#����@�����,b>l�0"OV�@%�v� ��ʆAYz�3�"O���Q��3�A8�� h]H�2�"O��`���_��t�U��)(�"OL�JǏ�E������׉Z�4�"O��BUo�@eL�5-r�ɩ"O���d0�F%��D��a�� �"OƩ���-Sn��'�5f�	3�"OX� ޞ6��)�&]���ը"O� ��d��*:B�)pƁ�J`Đ��"O���@%W=���+rd���5�F"O����/�7n���c��;yw�| �"O2x�C��_l)�ѧ��k�>��""O�)h@� ,ϰl���%L�ڡ��"ON�;�J#��9���\ȢL�t"O�;�&C_��3BJ߭C�4LR�"Oy���0R�!A�I���r�"O�t��ֿU��x��I^N2ع�"O��J�Ƀ�B�<}��읣R�`!�"O��ѣhC�gA�(+���9��RC"O��hc"Ԑw�6�V��K� �RC"O=�Q��36�+5��-���K"O.��� � �VyrV+K�w�2�8�"OFDr ��6-���$

�Vj���"Oh�5��,E(��CYP^�e�P"O�$ �ʔ4.8{���UF�y��"O�����<0Ys��'.$�(�"O�$�v_
;� � ��Kq�1�"O� � �gf�~�j�c�F\�Iz"OƸ� �-{s�cʖ0G�H"OJ���êW#<83ɔ(X#���"OJ�ڕ�L�T���rS�f�a�"O���e��)oY��c�|��!"O����G�g��	 uoL/ *@��"OB����C�j�|��0%��[��\i�"O���F��
7����΅2�"Ot=��lݛ)���aC)�h�x�"O8���тGsD"�P�<�V+V"O����[c����/!˨i�"O��!�[a�.����b��8&"Or VaWG�4��G�ɩ}SF�{�"OB��a,ۤ����+y���%"O���7�L�;U<����8���"OV��%
�T8pFʪ,��Q��"O�1`�7qk�ܪ����g"O��*�n4g� ��ЮP"��-�%"O�ȩ�B�5�8�Ɥk�̼"OhD)�n�	 xZ��ビ�ap�4"1"O�@saMT�)8��R�ȸ$O�a��"O���^2+�� P�J)h���"O����۪y��4�R���MztI�R"O�HRHπ4L���]� r~Xu"O�))$ �,n��ۨ4Ŵ��c"OzE8� ��7)&�8@"�$Ѵ��s"O�A"rɝ&K�H#�ǜ�)�V��"O���$ �:~��6��4� �"O��1`��S��	a*�p����2"OlxbL��Jt�� S�J{���7"O �Q��]*'�(!��/��`�-�a"O�<�� ɫ7���PAiQ9NLh��"OF9���ZdN�(���<P�Y��"Ox�����c�$�B�.���0�"Oj��p��4��2�F�7�4�"Oδs������Z��ݢj�^숷"O"��%ŊM��Ù^u|�['"OB!2[ :��y�Ȋ/"^p�(&"O:�S""��P�F�:HA�A�"O��1�`G3>,���M'F("D�"O�a�6)ֵ7�.#j֕څ�1"Ox�+dᓣ\,��8`W�rHA�"O����ɟ6C���B���z<�H�"O=�5$�5��h���.)�ȩ��"O�]���O40�\�y�	F�Dt�"O �8g�T4��	 Cʠ1xlɨ"O�����:[~QFL}l@Y"O2�R��sȡ�˂jNE��"O2 @���j&8�q˟�� h�"O���ą1I��� RD��k$"O�P��*۲s��q��E� :�F5�c"OH�3�4R_�]@����0R�͢�"O�<j�W�(g(�R�!N����"OPPBB��c��T�BK^E,d�G"O�h���xzg��?��t��"O�T"$�Z2�੃�J3(��	��"O:��S��|�ʴ�d�Nl�Fe�"O  *w�HJ�h�Q�E ���02"Or�
S���(0�e0i��Dj��*w"Ol���� ?Q�j�rCHR
�x��@"O��կD�uHR!1���� �X��W"O(�˰c�A�<�䅇0�b�H�"O�DR��ݖk<���`��#����Q"O�"D�P�pب!s��1�u�6"O� h�q��\,�0�W�ގF��Z�"O��'�Ѫi5b�qB��'�x�`�"Ot�I @Æ(L.ؐVe�-p��s�"OH��t���;  \�FZk4���"O:h"�aH���Q�i�V B@�"Op$f��B\e�Q��'y�\5�"O���h�ȝє圓8$��,�!�y"@�2p��C�ґ� %Ѷ�B��cI��r�F����[Ӏ�|-�C��!��(2�Ȭ:��ej¯�.�dC�I�~�TY:�k�n����E�4a�lB��rJNŲƕ2��i3#d�/EBB�ɯg���r"f�=1k�	R���B�>B䉡7��!��ɘ0P�p�ɶ��z8B�	/_�n�pg��-zT�2mX	H�C��=E}.TH�\,H��T�E�6h��C�	�WbN���$�,�q�gɺE�C�	��ԀCő~G���T6FɈC䉭ft%ݦq�n�0�hE�~@�C�ɿ@�%j.�WP��!R�C��3]�V����%��-���Z�C�ɤb�p(�e�дN����ݴ9�C�I�XS����A|�q��N�)i00B�=y��jF�#cZ��I��U�U��C�I2H��ZdCN8	
�]2�S�ٌC�	������G���W��zd�C�Ɂ<J�)@`J�19n���XO�C�I�~�����Q�B\�+�-w�bC�	�oN����SF
��6ĝ?}�$C�ɳ#��tBw	�>��RF r&�C�	�t��}�i��vڜ}���\�O��C�O+u���DHvjtƞ�+�dC��4u=
y0�N B�J%A@M�@�C��:"ֽ8����q�nTp��]�Cu�B�	0}^�ɦ@ #�`����� 4��B�I%Gl��!vK�	b}�`��6e��C�I�u�@�E�-=ȸK�Q;/[�C�I�'. �u�:��e8��Ϻ>A&C��5}"as2��#�j}ʍ#,�C�	-�Z����N]�L0s�B�	���)��	LjP���_�iv"C�I�'�pSaKU5$�|�vL�2)C�;"i�ЇFF��T�%�ڈC�Ό���킮X��l ���5	C�IV�R�j��ߝ-���"U(Q%I"�B�I?{.Z@��Ǐ}FT4�Ro���B�Ʉ�$=���nm�X�@�kQ�B��i���5a�}�OC{�@C�		}��%��4�n幅l��c�0C�	6&�B�j�	�'/�4��Π"ODB�.�
y��ԛXqΈbQE��6B��6c�f�y�	�<x5�gK�w� B�	�j*0j?/��5H�E�B�I�,�$�㗠JL.�k��-K�B�0`T��ѢMR�MD�)x��	r�@C��(E;j٩�䒺L/$k��P��B�	3[ IS�XQ*l�a��B�I-j�ڤ��jV��g	�!<UDB䉮D�
J��;C�99�C�	�Q�p5*�˖�&*������B�C�	�M6����_�.�wL֚�\C�	5.+� �$�-$�D
��n�<C�	]�xH@���8�7Β	gf.C��4B&���Ǐ#-)�F��7�jB�)� "�; �F�%(��4=v8m"!"O�xsG&�y�Ta�c¨�z�"OhP���L��h@P���~WV�� "O4����V��J7�?M:�͸u"O ϒ6w��9%�	u��� �"O��1!�G&�l���cX�THMp"O��B^����0c"sr����"Or(+�� �v�иa��ݡLYx��"O
��taEbr�q�*V�sdHI��"O��!X�aQ̭��'ݾ	1nģ4"O�YJv�͈3�誔��5|Ԑ""O�� �K�>ta+��gSh��ǋ@�<)��O�9*0D�ufBM�������f�<���[��M􆓿GH!XpC�g�<�!Jا!�~�Jb���v<���Hm�<�tjCynڑ���F4&)���S�<��J�L����?���Ă=D�h� )�4EǞ '߁Q�9фG;D��b�a�<0�L���$LQc��4D��g@P65��l�Sl:k?p���'D�$2�o�,��y����h�Tx�`�&D�Xe%��^��C(l�F �s8D������D�Yc�E�P� �5D�l(�g��9Y"�� {�ęU@�]�<Y��I�7�X��T$�O]��xC���<a��ؑ�F��U=o�0��Gy�<�G�FzQ���� �8&��YY�GTs�<��mثpC"�r��\/a�nEo�<��?[i@�*BnMa�̑���i�<�'�V=sNz�&�S\ �� v\��0=i�م{�X���&�

XRq9�fn�<Y7���x�Jz֭رcZ		��a؞ �=)���nLpЋ��4ud �0c��yrL>w�:��m��b_�͓����>aH�����n"�U��vc���G+D��{�\�h`1�Rl�	RJ���P�;��hO��;e�`���#�(h������r�C�I�t��ȴ��8HZI���G(���hO�>5����$,F��Ԥ�Xm20!�O�B�I U�b�2��#�*-J��Y�	:C�9'Z�tjۨg���ubY9r�C�2�P�:f�P@;`@��ܞysўH����¾z9��٦�
�W7�ۀ�2{�!�$V+?��$ F��s�
�������d�U�9̑>�c�0�ۡG�~��(鶎J?g��)��&φ�C�*�*&V\�Ȳc�^��T`�颟H����v�es�&
�fMdXb��&*> �'��p�=)�m�w���G��;�v!�D{X��C�_��V���؀z&�[m�fQ#��7D���u֥c}
����23%)�(D��Ȣ(���B����=J�0���)ړ�0<�g� t`pc����u��!QV�<��CK#i��݋��Q�U���p$n�<�e!E1w}�ej�%�Bc-i��s�<ْ%Q	c�܉��I��8M��	�k�D�>٦Z�l :Q��JH�Xc��v�^j�<)�ղwF9yF����o���O<���a����4`�%(�?&�x�ҕ7�S��yr
	VhI˥N� ��U��U��E�?���s���f�I�M.6���'�tMX�	/D�Piuc�8P�ͳWVp��U��M-?YÓ5��[��a@ǫO���Kw/6�4���|�=�4�R�B8oW.`2D��
���FyB�|�2iρ2�<@śawR\����f�<� ���WL�1�H@J���j�5��"Oƨ��7+Cv:�:?ђ�i0"OTHK���}����C�܄ʓ"O�<" I�d4D��wO4m��q[�<O�=�'�?����򤝒P6 �'�3wΆ�30k+]!�$�E���"�a��X�00@�'�ҭD{���'����_
 on0�΀Q��������>MtDXde��
�2��	[�w��Io�����n�
)�p���m�$Li+8ړ�~b]��$>���C�8m�4A��	ZD���74������0J�L�b/��t6,h�c��f�D1�S�'40��,�������R����ȓ!d�y���0��� �kE�{!��)������!)>�Z�f��S��U�F8D���v�S�EPҁ�!��`��;�<9��F�s��YE��T�A@xĄ�yAP�H�@��h��^	N��ȓ\�*T�ĎF%J���I�jst($��D{��ti�
8�H�{�"?V�4�.Z
�y�O�73�H9��hP* x�)�������'|�zB���䨡0��Ig�ze90ʕ���=��{"��6 ޘ���D�*Z�xQ����yCv�څ��,Ŵ>�B w�@���?�'�80����=l��刣�f�D��	�'Ծ����0)*P�"˜�\��\��}��'�-��'�th<hSBlN�[���z	�'��y�����|�!-/%&�)��'��sa�ݕ/�`m��Ü�%�<Y��'��d�c6R,q4��2	��
�'.u*v!�z:���m�'>l��	�'�"���^�_�x�B#^?$DV�
�'��u�#�+|�4�#%��B��OB�=E��J�52��k�.�^y�e ���ybGY�(�l-Q!�W�0Dj�����D���DQ �p����;-���i�GA�a��\��tB��m e2���0|��<D�Pæ !G�&��Q�K�VX���b�>�7I1�O�<�c��p��[4+��yD��"O�+��\�d�"Xp N�X>ʈ�"O4�$�}p���U�e#���c"O�ѣW��� ��MF���xP"OM�(S&\,� ��޹1 Tä"O���%10��=ц��7-,�Jr"Of�fꈗ�.p9�+Y�xM	�"O`T#D��Ze�qY�@Q�8p"Op�4D�.?�jaq(ĸy�*�
a"O�11��7lM�D[�A�}prTc�"O>�鄠A �Ƅ2ᆎBf��S_�|��I<%k��˓��"P�͂j���C�7A�`���X�&,��2�l�&^�C��8x0XL��i)XqmI�a&�<t"O�|�f/�R�|p+�L7��<Z�Ob��;ct�Ӧ �@��b6aʫ�!�5W�pH&"^~����I��x�'Yʘ'A��Hw����*Q;���"5�y���<5�(%��;}���B�p<�N<	*O�T�e�R�<��F�08jZ"O���F�S95����fmE�"h�c�x�ȑ\���O�^��s;U�esq��7<�B�`�'i(�*4k�8�HK�ݟ8|-��4�hO?7-�>�h��]�Fn�Q�¤�%
�!��ң?�P��زf`H��L7%���Jy��'4�J%*TI�E�oG�U��|K�'�R���.:����5�ԫ}��ɒ�7D�� h�7o���.xb�]@2U��"O"�s�+�r��t���P?sU���c"O�pCR822%��Yl��W��kX�q!���A����GA?* ���E�;D����k��s<q��������x�È+K>���	R�p)!�A@��y�JƟyzt#�jޜv�E��m&�y� ��K�d�B�ᘂc�� C"���O(��M{��iгl8��#�@*� pVJ�0!��V�B��q¬��S�T� �A�Q�	]���xl1BSOM���W I�7k�s�"Oh�Zr�A)f����\6K�\�"O8���ݹXj��F؛rb�q��"O*�z&Z%aJ��G~P�E`v"O�8h4a�8F#t%s����x�@骥��.�S��>Xp�eـ�ѻ� ���LB�IW��D��B�) �<QB"=Q	�G�*]��S�B8����W� �`ц�vU�x����:�TTP��L:�X���$����A�7z+�4 �-G �`$�ȓp4����չj�|�rj�>_QQ��L�N`x��3id�5�B�~i�����T�?�T�!"^�st�9���s����K>��
G��T�qt�V2�B�N>�/O?�	�O%$��`��4Z�!e4��B�I�{������7���� Z>k�PB�ɕ"����5��?騜p����o(�B�I(o���c�D��	�W�ѵJ`�B��x=��I�쩇a�tB�	'7�,��E�Ky�MVB i�HB�I?6V�IA�C�Z�ĭ��^5�pC�	�|l�q�&F\�M������ j�B�	�M�6$Z��E�U�Zm��@�J��C�I�K�|8�c�hW`��Qn��T=`B�I�1I�Y��T0���8���(#C��5I[���qH؅%Բ��hߛp$�B�J�a ���e���p f� [5�B�Ɉ.G��Y�\�f7t�����2�B�	^�"D�F	�qP�}���H"o��B�	���a�%�#q��p���^NzB�� �Lh��o�
�R�;NK�1GlB�I�[��my�	<��(�S�	7V��B�I5����P�_�noh0�DJS;~g�B�ɜP(�����H
jLX�j�(�&�(C��%)�����V*�2�+�K�R�C�"i��H�r.,�h4����'X��C�	�i�����3)�
�FB��C�$�ڽ)u��X֐����O��C��&=��'�?�~��aB�i��C�1���5<
`튳o8~��B�I�ˆ���)�a�T�k�&�;5�B�I�J��,h@���Rݘ4�� [�B䉷|����|U�}���%.�B�&^
��j�O-Ef�����7h�C�	�s�-YUC�`	|�P�-6��C�	�d��-��%�6z�|�t.о
��B䉶w(�[f�ʰLz4�b#N��C�	I�vT�g.	/)v��,�1j�c��pR��m���􌆆y�,�b�&�I9���Rb��Q�@<8#��0eB��	
+"Y;_",lP�A
6xϪx�W"O@��2m�&ML�����;J �Ͳ"Oq3d��<TЅ��ڃMk��"O�� ��^�]�*<X�	3DX$"O�M����s�Z\�"^h윙"O� n��F�e�\��a�8ot��"O|�(�D�e�Xp��+��t*s"O�C-&l����ނs1�I�"O���X�|���_�Q[l�H�"ON�xg�ԫ�fUx!�P���"O��㱴�g��&�lw\yz"O��f�6<^a&�O��4|0G"O��A�I�!>#�pNL�:��k�"OX��Z��]\.���͇<':)��m4B\����"���s1�0�����)X��hÁ3�( C�у:I���� ���P;���S�<���ȓQN�e�Ѻm�i��l��IQ��ȓP @���ݺwAR%�d/>`.���|3�Y�P"M����b�_�@�X�����A�]�K�&� ;6��ȓX&�;Tl	�$&} �2D��|�ȓ��bF!	� U�$�W��eBd̈́�\X
1f�F�Fy�I�.z2H��CT���+3�b��͉O�.h�ȓeJ���GM�"�D� ��"�6���*t�]w�u�pE 1bk(��f�<D��Ԣ ��R��#b�%,iT�;D����YÄ���g�!�i��$D��b��2J��G.X�����"D�H�7�M�j��9ӣD�G*���5D��J�Ǚ�Q�蛱m�M�����>D��k�k�<� ��B�&��I��?D���88\�x�A.yn�!Sh=D��[�ш&���c�ȗ!�>�B",D�[F��b��-
�j�![<I��J!D�������D��q����,���C�O=D�H�7.[-`E^X{��|R�=i��8D��pH�?#�M!��7�f�Kk9D�DY�ʀ�Q2��5��q{Hщ� D�L��-�������$H�YY��!D��ȳ�?g
�͡�"քM�����l*D�$��"\p��/��G�D9@��)D��IEd�^�n8B��	*J��$:D�D�aJH12ǅ�4@(�ڕ#;D���Egꥠ#�I3�B�8D�x�pk��S��Y�A��1-�[u�7D�X�gʥ`�o�~�̑U�7D�	��Q "AaՈ]&<�<)��O2�ǐW����D��<B�bG6'��	�6ga{�$X1�u���ҟL8@�
�0��27!�W'�0A�?D� �P�I70��ϟN��S�1�	�jp�53��Q�)4LF����#Z$��CS�� 0j��^ �yQ�a���g)��(�GX�4�}qP	4lYT�`�ޢ|�'� �s�$&��Y��BND�`X
�'� 1� '���BV�����E��2� �Z�^=���'w��1�c�]���cլ�83�~�	�Z���:��t3�ِ�iu��Rꁺ -��H!'Áy(9�	�'/�m+p��m�x��ɝ�FxI>��i^!1bY4(�'4 �2�O�j���
��4 �,�Rœ�q/ ���'7N���b�24Vj���֐}��9Aѣ�<h$�s#�)�b�G�ݐ0@��N~�G���y�c�D�8M��-ɭ"$&�aT��*��x��"-|V���Fȷ`� �.��̲e �+zX��R	�c�$�"P@�X�<��*f���&HP��)���S�a6ĵ`�+><O�=�6'��g9ܝX�k^*i�
y��@tf���Bӳ^�ȁ1F�jȱ1�O(<���<�������d�;�@a��'�n�k!�g��飱i��5�R�-y d�Qlv>�Aa]��mh���L��i�2D����^�	M��[��^����S��) ����k�Ĉ�d��[x 2���}��6Zz<
��=C��m(�*�2�`(p��DO�R0 \�#�(��	F�? �u8��ş{�b=P#/6C�˲-�QJZ���4��ƈx^��*	
=��z���j�<�'��\� ^�8������hy(ӓJJAp�bF5�>�I�2���!�Jh�3��92F�2��\ϟ��A�2�&M�S��,2���S&~7�̣��Ӥ,y���h�~?������]6�G���+a�(�Ӏ��R��+�!1J�2f�?9�&�ʹ�t-ۃ��^e�I�w*,(Ag�%7��r�!̿SgL��dI{�Vh(����Ё��(�v(N�kҵq(��1,��@2 U` ��*qJ�$��	�!�V���Z
S{�)Q R�k�c�,AQ��,h��,�\���P�Y
,������(M�,O���@�	 +|���"O�YX@�Ľ3��T{�NEW)�5*d�� D�+Ӯ��b�L�!U"Y�Di�Q�~*�h�ۼ3F£N�2�Γ�`P�
�J�<q��]���
w˟E��)⃒ s h��[(s����1���'48!`�[��� J@��Nhf8�����L����� LO���tŖ%^[��Z@K��� !D����䉂m[<������=�r�H�qX��࣠_�C��f��F�t�+6�:�I�D�`�K���<�+���!cr �H�	�~�4'�{``M0W���h\�E@]��y"HԄgՈQY��\�z"�]�S�Pe86�զ���Ct����.v�^� v�̓�� h�B�&MB7Q<��L����~���^ T�6�)#K&%��[�i����x��� 3����L�	�O���e�� ��=�&P�1O�`��pM�����j�Z�;�&�2a��{��d��BO2a��m����;�$��橖8J�M��F�z̢�����I="�%a���'8lA�b&aޥ:3Ʉp��D!���k��p�U�!�Oj�H�
�c�´A� G���V)Ӯ"���yU&��M���	 ��P�I�J�V��`ʹM�X�>��P��1���z	���OhZ�P�*/x�J)�@��?z^�ȃ�'���Rc�>1
m�PLA#A�|��'I��P蚅gzׄ�Rs�?�� �^O���`S�	�,�3�*D��
��O���3�܁t�4TX�K�,"����?��5(g��f�����'�l���/;� ����,M⡡	�&���X���1(���F6MV� 'H0gȐ@�C�='bt�$sca{r�U�Xׄm���:���!�@.��O
��w��(ٴ��C��^>L �Ua�+x��Y�F�Q�S�H��d\���e�"O�8{A��eG�k)�!pdl9&�'�.�x��:b��1:�g�`Ԭ$C1h�
dF�5�W�ğX&���%��'f/+F���y��޴C�\�`�@B��r���Z���md�D�#  0z �X,��(�� ���!扙C��+U��Fr�UP0.��b]��?�.O��R�`X�iD�"�� ��A�|��,גU�%Y���386qpdL@�(�v���nzh��#��)X��|ʀ�ڲ<B�	���$�O�؁��9v��@�]�J>u;�ڟ)��4�7a�l�t�𫆖���GI��x��Mw��aYT	rY��?�D����dYpFE �&���X�'�K}�(W��i�I��=y�.4S#��]d�88�)lO�˓'M��D�
 Yj�r��*3�H��d�$]SЈ@��(bة:��E,?G�}��՟R9k@���M�K��W��,p.���'Q�l4�З2�I��MC�'�z�l6����R�xhh�ԃӣ�h�2DΘ=�N�٠lR$M6,
�� �*D����tӖ��$�<l#V���c�Ä5A�H΁(����O��'������b��H礆2eJ�1�#�
�.�,&{"��MT�2�d�I�U��7M/����B������"Ԏ.��<xS��O�q+ʊ*R͠r�4`����" ����˺��-���IܳpYp<H%#� m��3�&Öp�!�$��Mi��9d�
�D�}+f����Ԧ�ܟ�b$��a N����:���x�=�h��I���,���g���{"�'Ꚅ�EkO� �L�#�e��b��n���"�	�;A�o�p3��1'�xW�J�>X������O�*�D.Cx@
�A������'��8���gz� � ۅ>�VM�O�<��'w��9BRd/
��A%����s�O\ҁ㊚&s��7>B�D&>A�OC0XK�'�-E�zM�3,\n���'��e��ポ ��P���ێ!kE.X�7*�9pKy����X�����ZL�1����y���3iZ�]x�)�ȓx��-�!(Z���lz���vL�I2��EA/
'%a{" ��N�ZA˂��C�R(�
��p=�0��/W҅�gJˁ�M3 ��g����8�-S�ƛ��t��������_
bp��2��32J�&��3�i��x�jA�*l(�����O~��q�i���������'Y�P�'��1�6�6���2�#P/	hִ��\1m��S��^�S> 7-��v��kMZ�rl��^�지 ք�@[� �h�t#Z,�	2OԀ�`�2p>P�2��".J�iSS:`�T(��A�+����[?i�g�'!���6)�$hx8У�jR��1���V	;>@�$0s��Lc$�Z�p0��W\b�iA�~��Ƞ,�ڐb)tĻ�f��h�Q����J��@�'v��'E�T�H	 -+�#�92Ol�����8��+A#~�Zɂ�)
�&}Fz"�SzwQ?ecV*&	s0tq�Ȗ?Ք0�.D�dؐnX�c���fn�skR)pcl���C�O��	P?E��4���mB�y?��i�pv�Q�o�����I�;�t�óh�	o+�+�R�Z���ΓW�~�?�үU�!h6lI8KV�ч�[L�	�KWџ$���>�Z���PK�tJ"
�W��y��'�Ҋ��&~�!�N�m��2�G_X�J"=iUb�����x~B�i���0�R�;�H�B叕3��e[���0�'�L�Yb�;x�LX�w{�"P�'���,�Ms�����#�M`�(@.Л8��`�'�@�~�)B��??�ڷ1T�b0�Ԅ~�;c�X��yR�xb�rӀ�?	��Oc���-O<}P��U/��d;}��$*��صO��i��A�	�P����
O��7}��̹�l�o-���t�]!��Q�kӔc��̓e�D�d}Ӫե����X!W����	��f'��Qg�9��=af:�$Ǳ�JA���=.� �ↄ`8r�(���I
�yr�T?�d$k��Ի�؏}lY� ��,>�0h���?-��UL��鉤aA�sx�lKe'��d�=�Óe�,�C��.N�x#B˕5��[��)��P��&��w�6�h0LW)q��1IT�=D��P	�*��`ץYª�%�8D�,�c]�[��[0�X�\y!��2D���jF<`6���f�TKP�$k*D�XöBDd��y�J�8���k/D�h��aG��8�a�!W��q��*D����.!t츥@TbM[Lf�)�!/D��Ǳ'N��ЇQ#�6�Lw�<�S����pEo7 w�x!d�w�<��Ǚ%)�f�(��*��DW�<�-���E)���%B+������S}�
ax��"v)	;p���DڝʼԸ$�'�O�а4�g��YR�O+��9�g��r.�=
Å��\	6�'��Cw�\�}d�X��ăc�,|	��}��O���N�z0u���6p��hz�"O0�b�N"}� ��ւ,�5;�@#*g��(�'�>i��������	�j*�r�&�-,Ԏd9d��vB��B�<@$o��wb¦bH���C�	X�ZU�vjK��u`�`�l�bB�	3-�$ ��f�
8jI�(�saxB�I�v��{�U�&����dZ �ZB�I#2R��0��D�ȵ$�8�B�	#G`d���V�Z;J}�e�U�:��B䉇	h��!)z�(���L*>?�C���.���N�>�� ���{��C�I!Q���AV�(��a�잮�C�I�ب��"@5n�4j�(�2%�C䉕N�t�Z���}M�d袦��dC�IR�~�Z�j�7�=@���6�$C�ɇg�T� W�5F9#�Ʌ5�NB䉾g�`X�&�|�Kp��JC�I�3o(<�a+ە&��5WK �"B�ɉ`/r`%�	&eL���)X�Z�C䉢!�ȅ�lE6/D��V)V��C�	,�Yr��\ v$R`�A?��C�	-.�}P]���r�ĳ|�Ҡ#
�'O�uX�߁yH��V��_�5��'Y,1C�G΂4E�Շojȹ��� �X�1�:\��q"��6ܱ��"O�`r���@ܬ+"�	��E�W"ON!�6E2X�	G��"�;�"O��S�'ԶJ/n���&��Zv�!�"O���c�:L ���;V���"O��S�ː4wD��Պu5Ir"O��P�/��؋�B�<$�i�"O|U�g(��w> )Z�a�&��r"O2 ��#P�l�c@��~?.��"O���j�lɂ��E���"OD��r@�E�`�!���;�"O��P���"˹ՠȰ�hC�y"�-d�	��1эD+a��)[
�'��)�k��������$�`M@	�'�JV�	+�虨��- �p�'D�����D�J�X��#{z�H�" D�h���
��L	%B6 �.2%�;D�d��DƧp䐀�AR�TV^��@*D�8�S�η Dp�ۀ��/k�@�b�i)D�h�gN��������/TsLP���)D����IQ�i$��ϗ+��y��*D����)��HI e8JJ�ll	�S"?D�̸����ԅX�KR�HTi@E� D�4sE���&J�z �;]yH�brA;D��ś~�`��)V�f�Tt�gk,D��I�N�>~��eoB�pTL �d�(T���%�f�ڼr"7�}j�"O25ҶH� ����0�A  "O�t�T%ߜ�\l1'!�$$�&�[V"Oإ���t\0PaQ�Y�ZT�P"O����.>:�d8`cLi��� "Ox�8@$��,�Ty�v��)��T"OؽFO�.Y��;�kC�2��`�"O�v�X�H�E�!�� �����"O�k�gE�x~�,@� ~����"O��C�:9|p�&�A.#lh"O���`�T.1K��R��T44X�LɆ"O0��G�?�d���-)Z��"O&�`+X=8�>�Pբ�GB�j�"O��P�2S�Ț5��HA�"Ol�IV�ڕcNE�钟	}
��V"O��htJ�(T���2Ț�(4��"0"O2����3���/y?��A�ڋ�y�nۯ!�8� C�� 8����a��*�y�Nf��A�`��)+��Y�	�y2G�B3�h D锐
)�q�W�	�yr�ӭ��;t�Ń������yR%��ѴQ��A�s�����-N��?a0[d�\2�x|�9��M�A�&�5�N�p�4�퉄r�ȡ�N�g�OX �\�[E鈘r�,l���ș�yb �
A|uy��v3����mC0��'��q���؛ ��A��Ӆ;	4ea�ίR�Ƽ��C*
B��7uS��1%"�n8;���k��]���V:�1�(O��ˏ�Y�D��U�u�U��!d���4�<D��(�EK�.9<͛'!D=,q��*�F_�c\�\�RCҿL��
�R�H�q7.Nt�H� #"	U��q��I:u!N�q�	E)y�6���4J�����0���0�[)0�p���*H���VP2�e�P(�8�l�$�`� �J=�t��Q�C%hy�>Q�!W�3�Z{� � ��}+��6D�$R��I�%�
�2)�42�N$z!�� @�\	�m���~R�Q
���@B����� �a��E#.
���ƓsT��qύ�P�82��-���*���hjA�!1���X�RQh=�F�-3�q�פ
��ybb�,6�A��ԋ�����a~�h $\ w��QR�Q�0�!�� �Y:�ai]
5�q�2P$$J��|R�3U(<(*t�_$?����ۥCg"훱6!^��r*O����ɡy
�a�:Tc��9;P���P�X�0��B�g}��Cwp�@���D�Y��O¼6�D	#TG��	VL���!>*�bk�`�H�c�o��[Q������%��]8�Dx�%��IFI�4��!�-O�<;f�N�}'`�Iщj���"�'��4I�H4Ewr	� 	��xӍԠ\}�!
� '�E�'�bd��G)�n��FE B�Od�Tjr��6u�!��"_�� �{��։v���3�S:#t�	�\�4̙�V1Av�@` �0B���m�;�0�z"I�s��a�'����*�9�ܑ �'g�DzדwfTѐI�<�Z�c�ʟ2Z]��0�)֑S����ԅֵt�n�u%�U�l	)�e��`L^�8܃VO٠K�e�<�v�Y!H�}r�i��@��e�¾o���P?тq ý��pq�ܟ\	�$�*D�����e���҇�I�@Cҝ��l
�Xe�uq����~�k��\�mŸȍ�T�ڳ�yGO��e��c�B�$�5�����y�C�n�blU�Q�
wtU���0��&�ǅT-�0�W�/��`���ٌk�z"=)��ͦ�Q$�^?{�����ۍ�0=�O�G�R}����s�2� JT��T��Q�Ivz0�԰C�Hi3��1}Pa}B�_|AڳI Ǽ��ԁ�ܘ'Ŷؓ�Y��9�U�%?Κ� lK=M��3��	���*Wz�m��;.� C�	�U#xd�&�LQ���@��zT�
��Ɨ/b��iJ�{�6�^�O��Iћ'��]��H��; u�E��	P�'�zu�W�i4Lm��?N�Yy#��BH~����f8�|qqĈH�)�M{ ؛E)�<)�5/���	lP̫@��l}B,���F@��(��rWn�;�yQU,��f�� !�|����ۅ�ēA@v�2s�M7
�Z➜���E:�K�_�%�����,�h���e*H�/^P��6m�:�&�ʂiS5X�����o�!��-��D#p�H.EtD=��l�<Q���H�6=��rd�IF�=�@e[�7�\�Tk��%f!���fKڽ�RKW�N^raP�j߮?Q��UY�JD�2�ó��)ڧC�च���M�%I����@��!�ȓ2h� �0J�4M�1&�#=��OL}��1Ap&(9Óp4l
��5	n���`k�6,�(���(�*�p� �!�qboS1Jo�%��J�Y��1b�'�2���R؞L�lϪA�<�y"-�/ ���
 �<�/���J4�B�$��6픴_����Eٞ8$a���6����-&:�9�ȓgx��u@��T�~u�5�N^jD�� �b�K�,+t��Z�]0;�� @.�'x�,y�sw3bI@|�Մ�4w( 2���w\����ʛGcԱ@S�#��;�% h:��YfK�S��'I:����%ub%ʴ�,Y��Z�K>�Ã��d~D�
 �<�ʵ+�Z��D�+����ޫ�0=�ӂ�7�p� @^�#PR���
u8�Ha$�8,�����M�J�֍�Ƣ^�-{.�i����!���f�Ĝ���Y
QK� �ף�l�Q�(঩�`�Ѐ������G��|B�9�OD�s��C�	��b1�P�*]i�����3U�H�B�DxQN�6��S��?�D�־B�p0Ѓ3u �@��GF�<�Wn�T��Ѕ��i�
���h?��� �72Uw %LO*��Pm:����U�.�=;��'\ 4S&,W$w�r����B�� uŏ�P��- �M4D��WF� V��` ���&P?��q�>�{��A�5�'T���;T��|��A� ��m�$����2"Ο�w�ԋ��s��Y��:Yhm `��}��׈�&�~؆ȓ'ظ-��F08h�+�C^�g���6���Q��8�O�aSC��;ff���A�e#��{��'�
83�ޢf���V� ֮����%�R�+g ��y����8h0#ݧy�
e�@��.��'���5Ǔ�$%r%D��(W�G���y���rYl���$�yB�����Uk	=������A�`��)��]���'	�>�I#T��4�Ʈ�7Rʽ�ǌ��HtB�Ɏ~	�$"�6-��Yc�W�3W��$1C(Z\�B��4ǰ=Q�$��e^�e���ΰ*��@�w���Q�C,h�e{��� �]ct. 	/��Ur�,��5H�"O�5ذX�ػ��\�##��$Ģ ߺe�Q�H��y@�)Z�����p.47��"O�9x4B��F�Aag�
n�h�*�C)(�d��5�g?Q��:��tp�� 6��Y
U�d�< G܄��rT�N5���d�����,L0��'|�h��S�:��+�"�pY�\�e� K��?�7 �J�F�h6���|��I"�A'T����/J�0b,j��ǋ:�>�k��.�v[���*�i&��R(�|6*$i�/��x]J��ȓu�I����Vla1C�V!�y��K���A�� i\�å=�*���d;`ݫC/1z�JD�g!�u���ȓrV��[6 Ϫ]0) �/G��,��136p٦hǴ>R�|" �#"M�ȓ.���i���+�y��!�8����ȓ)��@�!&S9r����w!�/9����ȓ9XHy^8�m��*�$NZ$݆���ce��RHj�
��!Lb%��!�� ��>X�8DJȤ>2ژ��`�x��	X���.#G�A�ȓ?�� ¢	��:��L�uaG#t�lԇ���8JӁ��3J���b��W��ԇ�S>.-TC;A��j�I�*{���ȓN��<2�d��37����!(m�!�ȓ=����O(� 0W���Ex�ȓ`%V5���4l�`h��B!\�L�ȓ?��"R��0\j .�=�Ф�ȓkTP����n�h�w됟J,�фȓ���Z%& �<ڄ�%��Y.y��o��9ЃB�h�4��s�V�o����ȓEG�KE� 6��)e��c��U�ȓ7b�3D�B=m�nuib�;0޴x�ȓ>lP�ss�R9Ap��7i��ȓY���D<#��(�"�,����A`���%���9��$�Qƌ ��ȓIb�y愅1&<1��T�3����GF�)#D�ĔS���z6�+f��)��%D�Y�ǠJ�n�x��RF�
U������e�7�ױ_��zȧ�7��m��V�����1�����O8��@��n��p��Ǉr�8�cr	Y���ȓq5��ӂ(��V�\�S0D�-\���5K��`��>���K�MB�A��,�ȓ�J|ɓ/ӕmT|�Sh�F�h��}T
�i ��p�<�ȕ�؉5FE��\yx蠕@��dx�!��� JȄ�l�%;�D�o�>����͒`��#8pk��Y"�0�2#ʆ���m��yER<05l��KP\	�ĕ��=����Ѷ�J�9_�H�dg� z����r~p�q��i@i��])g'4q�ȓ]�4�@� X�\����nH�eS�Y��h�F�p	ŋ:����E)<*�$9��3G�D��.&H\�h��cI�4��'�	
P#J:8���
1S&F���mr� F��j��8����]bvp�ȓ$�����׋3��<C���z����YO�`#qC�?zx��r�:�ԇȓ|�Ys�O]vxY���U;6�
��ȓaJh� ��� Q@��#F �ȓ]�b0�C���;������5�8���@b�(1��ׄ��x`��߸5��ȓ9��xH�εT��(���9e�>���S�? 2թ3e�3���c�	�Zђ�Z$"O���эVf�)k$ Y
Bⲅ@$�䘉E�8�.���vI� ^1A1O5��D�w��y���j�B���"O� qO͌3^�H3�mT:%A�"O0)��Iѽ<,Rq�	�8j��G"O(X����j�p�1$>�	"O�q[1L�*5}�0�d֠}T�2F"O�(�f���5��iҤ$rF]��"Of�jF�`ݚՇ
=-o��9�"O��Ѭ+]��x��	@l�"OX�pDY�4T��v�ҭ"�D	�"O,$�D��Nr
���a�;<d([�"O�ݠ�`Ǆ_~�|�'�iV���CßM��z{j"|��O�\Y����|����L"1Z�$���E}��'i�O�$��21�J�s�Q>�������7�
�i	X�f�<a�o��+Y�!h�*_�y�GF}�O��b��M�3�r��dŐG�� �3A
�v��P2C�[LTq�� ɳ���� �\ ��
\X�h1'Ҽ+�h `n��@P�	�0|�SbԈ11n����H~� ��p�ق;$D���L}�F�����<|��8h��]
65��[G�P�����?OޡhC�H9u��1�?7�M�'\f�M�@J�	j�H��GӪX6Xe�u���T�T��>�T���
;�)Yt��=z�������3��RA[�P�6�N�t��c kEm>u��̟u=�q�˙(<Ԉ������Q�c^71����S�X�^N�����`t�T�Ջ:���dKO���YVg�_��ĩs��>�~
çA�y9eR4C�����۬qM0���CP$A;da���c��/�z=��G�C�!X`	 ��P�r��3^J~��'dx�.�H�S�JZ������*��Q�،L�0�z2V uY�4���-�M��I\&XNd��k��S��zW� "B�R�'o��;���'nG�,��"�`8q����5U>u3
�%)D�B�n(@�NC"|FP�ȓ}=F�0	4Cy�+�	�h指�%�t�r�fſ2p¤{5�.K�R9��>|IQ b� 
 ���  �df4�ȓ%��T�FĄ�ش:��G�,��ņ�!��A�S���zv�T��I/@P��ȓ�t�S!FZ=x�4�@��#�����U��!G�Ca:�!��D����h��ċ�� �@��ꀃX�L���"����w�81�0��	ɄZ<��<�Yi��	3U"Ҩ���Rv쵇ȓ}�!Aѐ^��ꆌ�D��!�ȓ2L��w-�Y+����/<1F���I#��I�(B,U���<�����Ra3�%M�jY�(� L9
�\��ȓi<�=BQiK dc�̓#�X-��݇ȓ	:���#?�ݑ%j,Z��Q��K H�(sj�(娙�O��ȓ9����O��t��3'�΄�Hه�ֺI��S{�!�5 �|�Q�ȓ��3n��v��P2�սY�X��U9δ#��0�
��QƆ<H�D1�ȓRCZ�K��/ĎM��ǴR�f8��r;���ɋ(Y ��b�'�1'�dل�,,)cUeS>JrlĂҫ�*��\�ȓE��p�&ED�� aL5�����y��ȹ�ۛ6c��
4-ʜQҥ��[tl��& ��(�����Kz���$Nhsqe��.<B���&D���)�0���Pu&ߍ���Qޠ�{W��>_<X�I� ݶ��ȓe�8�a�G��`�XR!��E�d���%��x��ݹz|��Y 2'��Q�ȓ1`�yXD����A�cݶQE�\��4>J�˕�M6�@�2n,E� �ȓ��!j��[�QoN�i5 ^�XY��R���I��vC^,���4Xd��S�? �$�Q�ez���%ꆞ���kf"O�re.T.��,������	��"OY(��qa�b/�{��@�	<D�4Yc��67T���&�� ����$%D� H���R� ��Ó�]� D��e=D����^�0����Ѝ-"�:Pn7D��G��1E�nq��)�/���2��4D��ypG9A��0��B�4�֌)!�3D�,����)~#��ypi 9=��肴a1D��Ŕ�}�d���ұx�h��4$D���✯}q:qq�E%rF�z��-D�X3�ƍ�$�"��7cΟ6��E�C0D�\J���o&`���˶L���c,0D�D��o��r߼t���Eid�@xF	#D���f	D��)�/P�����!D���5
Ηz���*��@(0:�ӗ�:D�dJ�L�D�!QfHx���6D�3��)d�,@I��-f�"ѯ*D��i$�Ę.twgJ�_�&ɱ�F)D��{���Hs�ɇ;��	p�+D��`@�+�4��F�D�"�@쀕�/D�p�Pc��y���voq��97'!D�H�R��+��Y	�E�C�剣�?D�d��	J p�����IR<~��˴�!D��+VbҧQn�ᇪL�W�F� :D�D9W �cPP��o@^���[�8D�4*�H�;�)1�/�#X�
�q�4D�@�p���c ꭱ+� Ac:�ð�4D��ȢGҖE�����c���$�c��4D�!KY�9x~��r��	��Y�f.D�$z�"�+Z;��*���h��8�q�-D�<�`��.B�����ƞ=e��@�7g,D��R�Ի�0��V�Ur�g'D�4���K2= }RLF�e�V 9�"#D��d�	o)�!�Į^�/c���*O���t�\�+�債��H*<A�6"O  �ƍ��g�l�����g��"O}��L�\������"OR�h3#� @��"f�4���"OؕJe�
6�AxF/�7`����"O^����-�p��	R'UFɕ"O
��e�DM�ݓa��K8���"O�I;�*ԝ]~
��m��78F�"O���#��dbH���,�X��(��"O�T;A��B����vLӚy�����"O�ٹU#S�$O��Ò˗�2��<Q`"O��7�Ϙ-�d��Rj��=����a"O�L�%n�13�I 1
@'����=�!�� �r�J�Y�*���<��aU��!�ۮb���q� We`���(UG�<9cb��1�B���JS3��M�E�E�<�@��`a+�gܙ!����<���em")R���'�hԛ$��y�<AAj�wE�\h2K� ҶjB��ȓ_.���j�V�@��U���Qʂ�ȓX,���Jޮ7i��
/��d��L�ȓzBh�R��ݫ!���W�A.5`T�ȓa�E���ɒ�U&)qB���ȓ,�N9�TļG,2|�ƭ'}n���8ZE�a˂�i�ޘC@�H&p�P�ȓF���j�;.uj s��!`���ȓa�!��*�A"�c	�a4݄�uD�4)�Y���l�E:=a�ȓ5e����\�	��dȴ/t@��S�? ��)��FNY"t��!V��bP8B"O���_9C&N�1�f�&e��qr"O��"�%
5)�
7*˥qIf���7D��a��e��ꇦH�yqo1D�L񖤖�s@<�s���HZ�p��"D��2Q׶b��$�! ¾x�
�{!;D�d7���)z.X�'ڈ��`���:D�Ap�@�RK����&��f:D�H��ɒM�TBϒ�O���k��6D� ��%Q�+�`�2,ϡ ����0D��bgE	.�2��TH�{������ D���B
${�0�!�L3uQ�tr��9D�(���4s����g؂9�(��/8D�X�uyI@����6@f�XUd5D���'f�+���x5jR�7\�P���2D�dywoC)nw(�w!�6gF�[�"+D� �Q��b+ p�%�Q��d�`�>D�$;w�Z�\� ��ajMI%z���=D��h�DB�|Ҍ!m�-vD�ذ��:D�p+EMݢq�����"O�̨�TG,D�8�d!�#I0��pՉN	c�v�2Di?D�$T��5ZN�Bm̺����T�1D�x����J�L���VUV]��/2D����͆$:�r)��LI��&4D���f֩U�rĳpgZ�mT U+f�0D��B���/'�#�e��Y̼ `N:D�6�G=�����b��K=���c#D� Y��@�0轺�-ͽI�ptL6D�8�ot4�� a�M�F(|��B6D�h)��
="-�l+�H
;��X�6D������4�ĀpU��Q��J�5D�X!á=mK�܉��i���{�e8D���j[�8'&?֖��(D��06�[1}*11C�?���g+D�8(SO���SnM1{�Z�*%�;D�,Q� T���9b,َsp�A�:D���ለ3U�t��늄*�l�x��6D�p�rD�)�\���H�wRXHҧ2D��{��wW>`H��H9�Z��.D�0� �}�Lq��DE�],� iPk.D�`�!�ո��䈕�ը'p��&7D��C�c��G�HӁ��wN@��"D�<�bO�R�&��0�Ιi�P�b D��𲈞�{�R����*|�ر�a�+D�`�+B��
��u�Z��I+�'D��� b���^$�!`��4a"D�L+ �@��6!��@�Dt�
��:D��)'��$�B-��G^<4��E���7D���UƝ3 ��=�&��?0�\Q⦄5D��x��ʰ��
Po��).����5D�\׈�"�� `cM�2�,(f7D���A�ʛ; !�N�"4�La�	6D�$
��^?-m�x� k�����,2D���DV�~R6�G�;"�Y��+D����j6<�<5��O�88�m�U�6D�d"�'R�E� !������)D�T�#eԳ�X@{fS�h8���1D�\�a�h3���G+��i�Rl�V�;D�\�РM�[��88Ga��(+@@���;D���®�F���1D�:l� �b�.D��y׊��0�Wq���/D�Ha1�I'G�J9���Z�� �!D�
�g��~��32��-z�!D�t1�[.cyP�H#gV�q�l���A;D�� �M��Q�u��uqk_'NJ�t!"OJ؋��\�b�@9�#pC�c"O~�r�F�8�Ĩ�t��L�L	1�"O��ZC�1	+�)��MV�P[��ڶ"Oj,�(��U\�*�8*dYP@"O�j��A�;���q.�:b"O�(��JQ'�N #Q'[`�@�A"O��K.�w"�0j��J�l�,Z�"O|L��D����� M�1S��� �"O"4
�\�a1�yAk�2R�)h"O�:D͖(A�^���V�A�Y�t"O���<r��E�&Jf��	�"O�\j灛�nY�(y��R�Zh� �"OZ)8�n�7$P�qr"�C��`"O�QY ��!'$@��T��wڲ�q"OJ�u B�tf�9��'"q�2�"Ov�Y��Y���`�K#bn2�3"O����[�$�1����|�����"O�U��χ�&��q�m� on��%"O��Ȃ7�M#�.��F��mӱ"O���!��;�,Y4�Q����"O�I
��Y~Z	Sヿ>��@3�"O	�NĊQ���QÌ̽R��1��"O� ���l���L�P|�y2"O���9�(� ��9��b'"O�C���	�L���\�`�L�J�"O�ę��J�L�`DE<D����"O�"d���Ru�ڨ;����+D��R&E[3j֍H��E�d��xRA�?D�x�@�;0��e�D�r7�3�N9D�\�U��E����wM���완�<D�d��   �